   
    parameter PROC_NUM = 35;
    parameter ST_IDLE = 2'b0;
    parameter ST_DL_DETECTED = 2'b1;
    parameter ST_DL_REPORT = 2'b10;
   

    reg find_df_deadlock = 0;
    reg [1:0] CS_fsm;
    reg [1:0] NS_fsm;
    reg [PROC_NUM - 1:0] dl_detect_reg;
    reg [PROC_NUM - 1:0] dl_done_reg;
    reg [PROC_NUM - 1:0] origin_reg;
    reg [PROC_NUM - 1:0] dl_in_vec_reg;
    integer i;
    integer fp;

    // FSM State machine
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            CS_fsm <= ST_IDLE;
        end
        else begin
            CS_fsm <= NS_fsm;
        end
    end
    always @ (CS_fsm or dl_in_vec or dl_detect_reg or dl_done_reg or dl_in_vec or origin_reg) begin
        NS_fsm = CS_fsm;
        case (CS_fsm)
            ST_IDLE : begin
                if (|dl_in_vec) begin
                    NS_fsm = ST_DL_DETECTED;
                end
            end
            ST_DL_DETECTED: begin
                // has unreported deadlock cycle
                if (dl_detect_reg != dl_done_reg) begin
                    NS_fsm = ST_DL_REPORT;
                end
            end
            ST_DL_REPORT: begin
                if (|(dl_in_vec & origin_reg)) begin
                    NS_fsm = ST_DL_DETECTED;
                end
            end
        endcase
    end

    // dl_detect_reg record the procs that first detect deadlock
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            dl_detect_reg <= 'b0;
        end
        else begin
            if (CS_fsm == ST_IDLE) begin
                dl_detect_reg <= dl_in_vec;
            end
        end
    end

    // dl_detect_out keeps in high after deadlock detected
    assign dl_detect_out = |dl_detect_reg;

    // dl_done_reg record the cycles has been reported
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            dl_done_reg <= 'b0;
        end
        else begin
            if ((CS_fsm == ST_DL_REPORT) && (|(dl_in_vec & dl_detect_reg) == 'b1)) begin
                dl_done_reg <= dl_done_reg | dl_in_vec;
            end
        end
    end

    // clear token once a cycle is done
    assign token_clear = (CS_fsm == ST_DL_REPORT) ? ((|(dl_in_vec & origin_reg)) ? 'b1 : 'b0) : 'b0;

    // origin_reg record the current cycle start id
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            origin_reg <= 'b0;
        end
        else begin
            if (CS_fsm == ST_DL_DETECTED) begin
                origin_reg <= origin;
            end
        end
    end
   
    // origin will be valid for only one cycle
    always @ (CS_fsm or dl_detect_reg or dl_done_reg) begin
        if (CS_fsm == ST_DL_DETECTED) begin
            for (i = 0; i < PROC_NUM; i = i + 1) begin
                if (dl_detect_reg[i] & ~dl_done_reg[i] & ~(|origin)) begin
                    origin = 'b1 << i;
                end
            end
        end
        else begin
            origin = 'b0;
        end
    end
    
    // dl_in_vec_reg record the current cycle dl_in_vec
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            dl_in_vec_reg <= 'b0;
        end
        else begin
            if (CS_fsm == ST_DL_DETECTED) begin
                dl_in_vec_reg <= origin;
            end
            else if (CS_fsm == ST_DL_REPORT) begin
                dl_in_vec_reg <= dl_in_vec;
            end
        end
    end
    
    // get the first valid proc index in dl vector
    function integer proc_index(input [PROC_NUM - 1:0] dl_vec);
        begin
            proc_index = 0;
            for (i = 0; i < PROC_NUM; i = i + 1) begin
                if (dl_vec[i]) begin
                    proc_index = i;
                end
            end
        end
    endfunction

    // get the proc path based on dl vector
    function [360:0] proc_path(input [PROC_NUM - 1:0] dl_vec);
        integer index;
        begin
            index = proc_index(dl_vec);
            case (index)
                0 : begin
                    proc_path = "kernel_pr_kernel_pr.kernel_pr_entry98_U0";
                end
                1 : begin
                    proc_path = "kernel_pr_kernel_pr.load_bipedge30_U0";
                end
                2 : begin
                    proc_path = "kernel_pr_kernel_pr.load_bipedge31_U0";
                end
                3 : begin
                    proc_path = "kernel_pr_kernel_pr.load_value32_U0";
                end
                4 : begin
                    proc_path = "kernel_pr_kernel_pr.load_value33_U0";
                end
                5 : begin
                    proc_path = "kernel_pr_kernel_pr.load_value34_U0";
                end
                6 : begin
                    proc_path = "kernel_pr_kernel_pr.load_value35_U0";
                end
                7 : begin
                    proc_path = "kernel_pr_kernel_pr.load_value36_U0";
                end
                8 : begin
                    proc_path = "kernel_pr_kernel_pr.load_value37_U0";
                end
                9 : begin
                    proc_path = "kernel_pr_kernel_pr.load_value38_U0";
                end
                10 : begin
                    proc_path = "kernel_pr_kernel_pr.load_value39_U0";
                end
                11 : begin
                    proc_path = "kernel_pr_kernel_pr.load_value40_U0";
                end
                12 : begin
                    proc_path = "kernel_pr_kernel_pr.load_value41_U0";
                end
                13 : begin
                    proc_path = "kernel_pr_kernel_pr.load_value42_U0";
                end
                14 : begin
                    proc_path = "kernel_pr_kernel_pr.load_value43_U0";
                end
                15 : begin
                    proc_path = "kernel_pr_kernel_pr.load_value44_U0";
                end
                16 : begin
                    proc_path = "kernel_pr_kernel_pr.load_value45_U0";
                end
                17 : begin
                    proc_path = "kernel_pr_kernel_pr.load_value46_U0";
                end
                18 : begin
                    proc_path = "kernel_pr_kernel_pr.load_value47_U0";
                end
                19 : begin
                    proc_path = "kernel_pr_kernel_pr.write_back48_U0";
                end
                20 : begin
                    proc_path = "kernel_pr_kernel_pr.write_back49_U0";
                end
                21 : begin
                    proc_path = "kernel_pr_kernel_pr.write_back50_U0";
                end
                22 : begin
                    proc_path = "kernel_pr_kernel_pr.write_back51_U0";
                end
                23 : begin
                    proc_path = "kernel_pr_kernel_pr.write_back52_U0";
                end
                24 : begin
                    proc_path = "kernel_pr_kernel_pr.write_back53_U0";
                end
                25 : begin
                    proc_path = "kernel_pr_kernel_pr.write_back54_U0";
                end
                26 : begin
                    proc_path = "kernel_pr_kernel_pr.write_back55_U0";
                end
                27 : begin
                    proc_path = "kernel_pr_kernel_pr.write_back56_U0";
                end
                28 : begin
                    proc_path = "kernel_pr_kernel_pr.write_back57_U0";
                end
                29 : begin
                    proc_path = "kernel_pr_kernel_pr.write_back58_U0";
                end
                30 : begin
                    proc_path = "kernel_pr_kernel_pr.write_back59_U0";
                end
                31 : begin
                    proc_path = "kernel_pr_kernel_pr.write_back60_U0";
                end
                32 : begin
                    proc_path = "kernel_pr_kernel_pr.write_back61_U0";
                end
                33 : begin
                    proc_path = "kernel_pr_kernel_pr.write_back62_U0";
                end
                34 : begin
                    proc_path = "kernel_pr_kernel_pr.write_back63_U0";
                end
                default : begin
                    proc_path = "unknown";
                end
            endcase
        end
    endfunction

    // print the headlines of deadlock detection
    task print_dl_head;
        begin
            $display("\n//////////////////////////////////////////////////////////////////////////////");
            $display("// ERROR!!! DEADLOCK DETECTED at %0t ns! SIMULATION WILL BE STOPPED! //", $time);
            $display("//////////////////////////////////////////////////////////////////////////////");
            fp = $fopen("deadlock_db.dat", "w");
        end
    endtask

    // print the start of a cycle
    task print_cycle_start(input reg [360:0] proc_path, input integer cycle_id);
        begin
            $display("/////////////////////////");
            $display("// Dependence cycle %0d:", cycle_id);
            $display("// (1): Process: %0s", proc_path);
            $fdisplay(fp, "Dependence_Cycle_ID %0d", cycle_id);
            $fdisplay(fp, "Dependence_Process_ID 1");
            $fdisplay(fp, "Dependence_Process_path %0s", proc_path);
        end
    endtask

    // print the end of deadlock detection
    task print_dl_end(input integer num, input integer record_time);
        begin
            $display("////////////////////////////////////////////////////////////////////////");
            $display("// Totally %0d cycles detected!", num);
            $display("////////////////////////////////////////////////////////////////////////");
            $display("// ERROR!!! DEADLOCK DETECTED at %0t ns! SIMULATION WILL BE STOPPED! //", record_time);
            $display("//////////////////////////////////////////////////////////////////////////////");
            $fdisplay(fp, "Dependence_Cycle_Number %0d", num);
            $fclose(fp);
        end
    endtask

    // print one proc component in the cycle
    task print_cycle_proc_comp(input reg [360:0] proc_path, input integer cycle_comp_id);
        begin
            $display("// (%0d): Process: %0s", cycle_comp_id, proc_path);
            $fdisplay(fp, "Dependence_Process_ID %0d", cycle_comp_id);
            $fdisplay(fp, "Dependence_Process_path %0s", proc_path);
        end
    endtask

    // print one channel component in the cycle
    task print_cycle_chan_comp(input [PROC_NUM - 1:0] dl_vec1, input [PROC_NUM - 1:0] dl_vec2);
        reg [416:0] chan_path;
        integer index1;
        integer index2;
        begin
            index1 = proc_index(dl_vec1);
            index2 = proc_index(dl_vec2);
            case (index1)
                0 : begin
                    case(index2)
                    19: begin
                        if (~kernel_pr_entry98_U0.H_write0_out_blk_n) begin
                            if (~H_write0_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write0_c_U' written by process 'kernel_pr_kernel_pr.write_back48_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write0_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write0_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write0_c_U' read by process 'kernel_pr_kernel_pr.write_back48_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write0_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~kernel_pr_entry98_U0.hyperedge_size_out_blk_n) begin
                            if (~hyperedge_size_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c_U' written by process 'kernel_pr_kernel_pr.write_back48_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c_U' read by process 'kernel_pr_kernel_pr.write_back48_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back48_U0_U.if_full_n & kernel_pr_entry98_U0.ap_start & ~kernel_pr_entry98_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_write_back48_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back48_U0_U' read by process 'kernel_pr_kernel_pr.write_back48_U0',");
                        end
                    end
                    20: begin
                        if (~kernel_pr_entry98_U0.H_write1_out_blk_n) begin
                            if (~H_write1_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write1_c_U' written by process 'kernel_pr_kernel_pr.write_back49_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write1_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write1_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write1_c_U' read by process 'kernel_pr_kernel_pr.write_back49_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write1_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~kernel_pr_entry98_U0.hyperedge_size_out1_blk_n) begin
                            if (~hyperedge_size_c850_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c850_U' written by process 'kernel_pr_kernel_pr.write_back49_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c850_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c850_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c850_U' read by process 'kernel_pr_kernel_pr.write_back49_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c850_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back49_U0_U.if_full_n & kernel_pr_entry98_U0.ap_start & ~kernel_pr_entry98_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_write_back49_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back49_U0_U' read by process 'kernel_pr_kernel_pr.write_back49_U0',");
                        end
                    end
                    21: begin
                        if (~kernel_pr_entry98_U0.H_write2_out_blk_n) begin
                            if (~H_write2_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write2_c_U' written by process 'kernel_pr_kernel_pr.write_back50_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write2_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write2_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write2_c_U' read by process 'kernel_pr_kernel_pr.write_back50_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write2_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~kernel_pr_entry98_U0.hyperedge_size_out2_blk_n) begin
                            if (~hyperedge_size_c851_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c851_U' written by process 'kernel_pr_kernel_pr.write_back50_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c851_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c851_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c851_U' read by process 'kernel_pr_kernel_pr.write_back50_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c851_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back50_U0_U.if_full_n & kernel_pr_entry98_U0.ap_start & ~kernel_pr_entry98_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_write_back50_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back50_U0_U' read by process 'kernel_pr_kernel_pr.write_back50_U0',");
                        end
                    end
                    22: begin
                        if (~kernel_pr_entry98_U0.H_write3_out_blk_n) begin
                            if (~H_write3_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write3_c_U' written by process 'kernel_pr_kernel_pr.write_back51_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write3_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write3_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write3_c_U' read by process 'kernel_pr_kernel_pr.write_back51_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write3_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~kernel_pr_entry98_U0.hyperedge_size_out3_blk_n) begin
                            if (~hyperedge_size_c852_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c852_U' written by process 'kernel_pr_kernel_pr.write_back51_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c852_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c852_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c852_U' read by process 'kernel_pr_kernel_pr.write_back51_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c852_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back51_U0_U.if_full_n & kernel_pr_entry98_U0.ap_start & ~kernel_pr_entry98_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_write_back51_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back51_U0_U' read by process 'kernel_pr_kernel_pr.write_back51_U0',");
                        end
                    end
                    23: begin
                        if (~kernel_pr_entry98_U0.H_write4_out_blk_n) begin
                            if (~H_write4_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write4_c_U' written by process 'kernel_pr_kernel_pr.write_back52_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write4_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write4_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write4_c_U' read by process 'kernel_pr_kernel_pr.write_back52_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write4_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~kernel_pr_entry98_U0.hyperedge_size_out4_blk_n) begin
                            if (~hyperedge_size_c853_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c853_U' written by process 'kernel_pr_kernel_pr.write_back52_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c853_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c853_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c853_U' read by process 'kernel_pr_kernel_pr.write_back52_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c853_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back52_U0_U.if_full_n & kernel_pr_entry98_U0.ap_start & ~kernel_pr_entry98_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_write_back52_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back52_U0_U' read by process 'kernel_pr_kernel_pr.write_back52_U0',");
                        end
                    end
                    24: begin
                        if (~kernel_pr_entry98_U0.H_write5_out_blk_n) begin
                            if (~H_write5_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write5_c_U' written by process 'kernel_pr_kernel_pr.write_back53_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write5_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write5_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write5_c_U' read by process 'kernel_pr_kernel_pr.write_back53_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write5_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~kernel_pr_entry98_U0.hyperedge_size_out5_blk_n) begin
                            if (~hyperedge_size_c854_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c854_U' written by process 'kernel_pr_kernel_pr.write_back53_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c854_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c854_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c854_U' read by process 'kernel_pr_kernel_pr.write_back53_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c854_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back53_U0_U.if_full_n & kernel_pr_entry98_U0.ap_start & ~kernel_pr_entry98_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_write_back53_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back53_U0_U' read by process 'kernel_pr_kernel_pr.write_back53_U0',");
                        end
                    end
                    25: begin
                        if (~kernel_pr_entry98_U0.H_write6_out_blk_n) begin
                            if (~H_write6_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write6_c_U' written by process 'kernel_pr_kernel_pr.write_back54_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write6_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write6_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write6_c_U' read by process 'kernel_pr_kernel_pr.write_back54_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write6_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~kernel_pr_entry98_U0.hyperedge_size_out6_blk_n) begin
                            if (~hyperedge_size_c855_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c855_U' written by process 'kernel_pr_kernel_pr.write_back54_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c855_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c855_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c855_U' read by process 'kernel_pr_kernel_pr.write_back54_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c855_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back54_U0_U.if_full_n & kernel_pr_entry98_U0.ap_start & ~kernel_pr_entry98_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_write_back54_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back54_U0_U' read by process 'kernel_pr_kernel_pr.write_back54_U0',");
                        end
                    end
                    26: begin
                        if (~kernel_pr_entry98_U0.H_write7_out_blk_n) begin
                            if (~H_write7_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write7_c_U' written by process 'kernel_pr_kernel_pr.write_back55_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write7_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write7_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write7_c_U' read by process 'kernel_pr_kernel_pr.write_back55_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write7_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~kernel_pr_entry98_U0.hyperedge_size_out7_blk_n) begin
                            if (~hyperedge_size_c856_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c856_U' written by process 'kernel_pr_kernel_pr.write_back55_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c856_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c856_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c856_U' read by process 'kernel_pr_kernel_pr.write_back55_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c856_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back55_U0_U.if_full_n & kernel_pr_entry98_U0.ap_start & ~kernel_pr_entry98_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_write_back55_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back55_U0_U' read by process 'kernel_pr_kernel_pr.write_back55_U0',");
                        end
                    end
                    27: begin
                        if (~kernel_pr_entry98_U0.H_write8_out_blk_n) begin
                            if (~H_write8_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write8_c_U' written by process 'kernel_pr_kernel_pr.write_back56_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write8_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write8_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write8_c_U' read by process 'kernel_pr_kernel_pr.write_back56_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write8_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~kernel_pr_entry98_U0.hyperedge_size_out8_blk_n) begin
                            if (~hyperedge_size_c857_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c857_U' written by process 'kernel_pr_kernel_pr.write_back56_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c857_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c857_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c857_U' read by process 'kernel_pr_kernel_pr.write_back56_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c857_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back56_U0_U.if_full_n & kernel_pr_entry98_U0.ap_start & ~kernel_pr_entry98_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_write_back56_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back56_U0_U' read by process 'kernel_pr_kernel_pr.write_back56_U0',");
                        end
                    end
                    28: begin
                        if (~kernel_pr_entry98_U0.H_write9_out_blk_n) begin
                            if (~H_write9_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write9_c_U' written by process 'kernel_pr_kernel_pr.write_back57_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write9_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write9_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write9_c_U' read by process 'kernel_pr_kernel_pr.write_back57_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write9_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~kernel_pr_entry98_U0.hyperedge_size_out9_blk_n) begin
                            if (~hyperedge_size_c858_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c858_U' written by process 'kernel_pr_kernel_pr.write_back57_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c858_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c858_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c858_U' read by process 'kernel_pr_kernel_pr.write_back57_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c858_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back57_U0_U.if_full_n & kernel_pr_entry98_U0.ap_start & ~kernel_pr_entry98_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_write_back57_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back57_U0_U' read by process 'kernel_pr_kernel_pr.write_back57_U0',");
                        end
                    end
                    29: begin
                        if (~kernel_pr_entry98_U0.H_write10_out_blk_n) begin
                            if (~H_write10_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write10_c_U' written by process 'kernel_pr_kernel_pr.write_back58_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write10_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write10_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write10_c_U' read by process 'kernel_pr_kernel_pr.write_back58_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write10_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~kernel_pr_entry98_U0.hyperedge_size_out10_blk_n) begin
                            if (~hyperedge_size_c859_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c859_U' written by process 'kernel_pr_kernel_pr.write_back58_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c859_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c859_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c859_U' read by process 'kernel_pr_kernel_pr.write_back58_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c859_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back58_U0_U.if_full_n & kernel_pr_entry98_U0.ap_start & ~kernel_pr_entry98_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_write_back58_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back58_U0_U' read by process 'kernel_pr_kernel_pr.write_back58_U0',");
                        end
                    end
                    30: begin
                        if (~kernel_pr_entry98_U0.H_write11_out_blk_n) begin
                            if (~H_write11_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write11_c_U' written by process 'kernel_pr_kernel_pr.write_back59_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write11_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write11_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write11_c_U' read by process 'kernel_pr_kernel_pr.write_back59_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write11_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~kernel_pr_entry98_U0.hyperedge_size_out11_blk_n) begin
                            if (~hyperedge_size_c860_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c860_U' written by process 'kernel_pr_kernel_pr.write_back59_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c860_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c860_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c860_U' read by process 'kernel_pr_kernel_pr.write_back59_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c860_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back59_U0_U.if_full_n & kernel_pr_entry98_U0.ap_start & ~kernel_pr_entry98_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_write_back59_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back59_U0_U' read by process 'kernel_pr_kernel_pr.write_back59_U0',");
                        end
                    end
                    31: begin
                        if (~kernel_pr_entry98_U0.H_write12_out_blk_n) begin
                            if (~H_write12_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write12_c_U' written by process 'kernel_pr_kernel_pr.write_back60_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write12_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write12_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write12_c_U' read by process 'kernel_pr_kernel_pr.write_back60_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write12_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~kernel_pr_entry98_U0.hyperedge_size_out12_blk_n) begin
                            if (~hyperedge_size_c861_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c861_U' written by process 'kernel_pr_kernel_pr.write_back60_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c861_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c861_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c861_U' read by process 'kernel_pr_kernel_pr.write_back60_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c861_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back60_U0_U.if_full_n & kernel_pr_entry98_U0.ap_start & ~kernel_pr_entry98_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_write_back60_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back60_U0_U' read by process 'kernel_pr_kernel_pr.write_back60_U0',");
                        end
                    end
                    32: begin
                        if (~kernel_pr_entry98_U0.H_write13_out_blk_n) begin
                            if (~H_write13_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write13_c_U' written by process 'kernel_pr_kernel_pr.write_back61_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write13_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write13_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write13_c_U' read by process 'kernel_pr_kernel_pr.write_back61_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write13_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~kernel_pr_entry98_U0.hyperedge_size_out13_blk_n) begin
                            if (~hyperedge_size_c862_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c862_U' written by process 'kernel_pr_kernel_pr.write_back61_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c862_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c862_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c862_U' read by process 'kernel_pr_kernel_pr.write_back61_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c862_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back61_U0_U.if_full_n & kernel_pr_entry98_U0.ap_start & ~kernel_pr_entry98_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_write_back61_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back61_U0_U' read by process 'kernel_pr_kernel_pr.write_back61_U0',");
                        end
                    end
                    33: begin
                        if (~kernel_pr_entry98_U0.H_write14_out_blk_n) begin
                            if (~H_write14_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write14_c_U' written by process 'kernel_pr_kernel_pr.write_back62_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write14_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write14_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write14_c_U' read by process 'kernel_pr_kernel_pr.write_back62_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write14_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~kernel_pr_entry98_U0.hyperedge_size_out14_blk_n) begin
                            if (~hyperedge_size_c863_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c863_U' written by process 'kernel_pr_kernel_pr.write_back62_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c863_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c863_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c863_U' read by process 'kernel_pr_kernel_pr.write_back62_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c863_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back62_U0_U.if_full_n & kernel_pr_entry98_U0.ap_start & ~kernel_pr_entry98_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_write_back62_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back62_U0_U' read by process 'kernel_pr_kernel_pr.write_back62_U0',");
                        end
                    end
                    34: begin
                        if (~kernel_pr_entry98_U0.H_write15_out_blk_n) begin
                            if (~H_write15_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write15_c_U' written by process 'kernel_pr_kernel_pr.write_back63_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write15_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write15_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write15_c_U' read by process 'kernel_pr_kernel_pr.write_back63_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write15_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~kernel_pr_entry98_U0.hyperedge_size_out15_blk_n) begin
                            if (~hyperedge_size_c864_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c864_U' written by process 'kernel_pr_kernel_pr.write_back63_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c864_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c864_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c864_U' read by process 'kernel_pr_kernel_pr.write_back63_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c864_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back63_U0_U.if_full_n & kernel_pr_entry98_U0.ap_start & ~kernel_pr_entry98_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_write_back63_U0_U.if_read) begin
                            $display("//      Blocked by full output start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back63_U0_U' read by process 'kernel_pr_kernel_pr.write_back63_U0',");
                        end
                    end
                    3: begin
                        if (~kernel_pr_entry98_U0.V_read0_out_blk_n) begin
                            if (~V_read0_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.V_read0_c_U' written by process 'kernel_pr_kernel_pr.load_value32_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read0_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~V_read0_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.V_read0_c_U' read by process 'kernel_pr_kernel_pr.load_value32_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read0_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_kernel_pr_entry98_U0_ap_ready & kernel_pr_entry98_U0.ap_idle & ~ap_sync_load_value32_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value32_U0'");
                        end
                    end
                    4: begin
                        if (~kernel_pr_entry98_U0.V_read1_out_blk_n) begin
                            if (~V_read1_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.V_read1_c_U' written by process 'kernel_pr_kernel_pr.load_value33_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read1_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~V_read1_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.V_read1_c_U' read by process 'kernel_pr_kernel_pr.load_value33_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read1_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_kernel_pr_entry98_U0_ap_ready & kernel_pr_entry98_U0.ap_idle & ~ap_sync_load_value33_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value33_U0'");
                        end
                    end
                    5: begin
                        if (~kernel_pr_entry98_U0.V_read2_out_blk_n) begin
                            if (~V_read2_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.V_read2_c_U' written by process 'kernel_pr_kernel_pr.load_value34_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read2_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~V_read2_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.V_read2_c_U' read by process 'kernel_pr_kernel_pr.load_value34_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read2_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_kernel_pr_entry98_U0_ap_ready & kernel_pr_entry98_U0.ap_idle & ~ap_sync_load_value34_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value34_U0'");
                        end
                    end
                    6: begin
                        if (~kernel_pr_entry98_U0.V_read3_out_blk_n) begin
                            if (~V_read3_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.V_read3_c_U' written by process 'kernel_pr_kernel_pr.load_value35_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read3_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~V_read3_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.V_read3_c_U' read by process 'kernel_pr_kernel_pr.load_value35_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read3_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_kernel_pr_entry98_U0_ap_ready & kernel_pr_entry98_U0.ap_idle & ~ap_sync_load_value35_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value35_U0'");
                        end
                    end
                    7: begin
                        if (~kernel_pr_entry98_U0.V_read4_out_blk_n) begin
                            if (~V_read4_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.V_read4_c_U' written by process 'kernel_pr_kernel_pr.load_value36_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read4_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~V_read4_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.V_read4_c_U' read by process 'kernel_pr_kernel_pr.load_value36_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read4_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_kernel_pr_entry98_U0_ap_ready & kernel_pr_entry98_U0.ap_idle & ~ap_sync_load_value36_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value36_U0'");
                        end
                    end
                    8: begin
                        if (~kernel_pr_entry98_U0.V_read5_out_blk_n) begin
                            if (~V_read5_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.V_read5_c_U' written by process 'kernel_pr_kernel_pr.load_value37_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read5_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~V_read5_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.V_read5_c_U' read by process 'kernel_pr_kernel_pr.load_value37_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read5_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_kernel_pr_entry98_U0_ap_ready & kernel_pr_entry98_U0.ap_idle & ~ap_sync_load_value37_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value37_U0'");
                        end
                    end
                    9: begin
                        if (~kernel_pr_entry98_U0.V_read6_out_blk_n) begin
                            if (~V_read6_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.V_read6_c_U' written by process 'kernel_pr_kernel_pr.load_value38_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read6_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~V_read6_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.V_read6_c_U' read by process 'kernel_pr_kernel_pr.load_value38_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read6_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_kernel_pr_entry98_U0_ap_ready & kernel_pr_entry98_U0.ap_idle & ~ap_sync_load_value38_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value38_U0'");
                        end
                    end
                    10: begin
                        if (~kernel_pr_entry98_U0.V_read7_out_blk_n) begin
                            if (~V_read7_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.V_read7_c_U' written by process 'kernel_pr_kernel_pr.load_value39_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read7_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~V_read7_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.V_read7_c_U' read by process 'kernel_pr_kernel_pr.load_value39_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read7_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_kernel_pr_entry98_U0_ap_ready & kernel_pr_entry98_U0.ap_idle & ~ap_sync_load_value39_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value39_U0'");
                        end
                    end
                    11: begin
                        if (~kernel_pr_entry98_U0.V_read8_out_blk_n) begin
                            if (~V_read8_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.V_read8_c_U' written by process 'kernel_pr_kernel_pr.load_value40_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read8_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~V_read8_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.V_read8_c_U' read by process 'kernel_pr_kernel_pr.load_value40_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read8_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_kernel_pr_entry98_U0_ap_ready & kernel_pr_entry98_U0.ap_idle & ~ap_sync_load_value40_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value40_U0'");
                        end
                    end
                    12: begin
                        if (~kernel_pr_entry98_U0.V_read9_out_blk_n) begin
                            if (~V_read9_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.V_read9_c_U' written by process 'kernel_pr_kernel_pr.load_value41_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read9_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~V_read9_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.V_read9_c_U' read by process 'kernel_pr_kernel_pr.load_value41_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read9_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_kernel_pr_entry98_U0_ap_ready & kernel_pr_entry98_U0.ap_idle & ~ap_sync_load_value41_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value41_U0'");
                        end
                    end
                    13: begin
                        if (~kernel_pr_entry98_U0.V_read10_out_blk_n) begin
                            if (~V_read10_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.V_read10_c_U' written by process 'kernel_pr_kernel_pr.load_value42_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read10_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~V_read10_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.V_read10_c_U' read by process 'kernel_pr_kernel_pr.load_value42_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read10_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_kernel_pr_entry98_U0_ap_ready & kernel_pr_entry98_U0.ap_idle & ~ap_sync_load_value42_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value42_U0'");
                        end
                    end
                    14: begin
                        if (~kernel_pr_entry98_U0.V_read11_out_blk_n) begin
                            if (~V_read11_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.V_read11_c_U' written by process 'kernel_pr_kernel_pr.load_value43_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read11_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~V_read11_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.V_read11_c_U' read by process 'kernel_pr_kernel_pr.load_value43_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read11_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_kernel_pr_entry98_U0_ap_ready & kernel_pr_entry98_U0.ap_idle & ~ap_sync_load_value43_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value43_U0'");
                        end
                    end
                    15: begin
                        if (~kernel_pr_entry98_U0.V_read12_out_blk_n) begin
                            if (~V_read12_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.V_read12_c_U' written by process 'kernel_pr_kernel_pr.load_value44_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read12_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~V_read12_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.V_read12_c_U' read by process 'kernel_pr_kernel_pr.load_value44_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read12_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_kernel_pr_entry98_U0_ap_ready & kernel_pr_entry98_U0.ap_idle & ~ap_sync_load_value44_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value44_U0'");
                        end
                    end
                    16: begin
                        if (~kernel_pr_entry98_U0.V_read13_out_blk_n) begin
                            if (~V_read13_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.V_read13_c_U' written by process 'kernel_pr_kernel_pr.load_value45_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read13_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~V_read13_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.V_read13_c_U' read by process 'kernel_pr_kernel_pr.load_value45_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read13_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_kernel_pr_entry98_U0_ap_ready & kernel_pr_entry98_U0.ap_idle & ~ap_sync_load_value45_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value45_U0'");
                        end
                    end
                    17: begin
                        if (~kernel_pr_entry98_U0.V_read14_out_blk_n) begin
                            if (~V_read14_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.V_read14_c_U' written by process 'kernel_pr_kernel_pr.load_value46_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read14_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~V_read14_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.V_read14_c_U' read by process 'kernel_pr_kernel_pr.load_value46_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read14_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_kernel_pr_entry98_U0_ap_ready & kernel_pr_entry98_U0.ap_idle & ~ap_sync_load_value46_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value46_U0'");
                        end
                    end
                    18: begin
                        if (~kernel_pr_entry98_U0.V_read15_out_blk_n) begin
                            if (~V_read15_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.V_read15_c_U' written by process 'kernel_pr_kernel_pr.load_value47_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read15_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~V_read15_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.V_read15_c_U' read by process 'kernel_pr_kernel_pr.load_value47_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read15_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_kernel_pr_entry98_U0_ap_ready & kernel_pr_entry98_U0.ap_idle & ~ap_sync_load_value47_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value47_U0'");
                        end
                    end
                    1: begin
                        if (~kernel_pr_entry98_U0.hv_bipedge_dram0_out_blk_n) begin
                            if (~hv_bipedge_dram0_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hv_bipedge_dram0_c_U' written by process 'kernel_pr_kernel_pr.load_bipedge30_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hv_bipedge_dram0_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hv_bipedge_dram0_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hv_bipedge_dram0_c_U' read by process 'kernel_pr_kernel_pr.load_bipedge30_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hv_bipedge_dram0_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~kernel_pr_entry98_U0.bipedge_size_out_blk_n) begin
                            if (~bipedge_size_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_size_c_U' written by process 'kernel_pr_kernel_pr.load_bipedge30_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_size_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_size_c_U' read by process 'kernel_pr_kernel_pr.load_bipedge30_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_kernel_pr_entry98_U0_ap_ready & kernel_pr_entry98_U0.ap_idle & ~ap_sync_load_bipedge30_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge30_U0'");
                        end
                    end
                    2: begin
                        if (~kernel_pr_entry98_U0.hv_bipedge_dram1_out_blk_n) begin
                            if (~hv_bipedge_dram1_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hv_bipedge_dram1_c_U' written by process 'kernel_pr_kernel_pr.load_bipedge31_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hv_bipedge_dram1_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hv_bipedge_dram1_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hv_bipedge_dram1_c_U' read by process 'kernel_pr_kernel_pr.load_bipedge31_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hv_bipedge_dram1_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~kernel_pr_entry98_U0.bipedge_size_out16_blk_n) begin
                            if (~bipedge_size_c865_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_size_c865_U' written by process 'kernel_pr_kernel_pr.load_bipedge31_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c865_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_size_c865_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_size_c865_U' read by process 'kernel_pr_kernel_pr.load_bipedge31_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c865_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_kernel_pr_entry98_U0_ap_ready & kernel_pr_entry98_U0.ap_idle & ~ap_sync_load_bipedge31_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge31_U0'");
                        end
                    end
                    endcase
                end
                1 : begin
                    case(index2)
                    0: begin
                        if (~load_bipedge30_U0.bipedge_blk_n) begin
                            if (~hv_bipedge_dram0_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hv_bipedge_dram0_c_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hv_bipedge_dram0_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hv_bipedge_dram0_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hv_bipedge_dram0_c_U' read by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hv_bipedge_dram0_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~load_bipedge30_U0.bipedge_size_blk_n) begin
                            if (~bipedge_size_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_size_c_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_size_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_size_c_U' read by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_bipedge30_U0_ap_ready & load_bipedge30_U0.ap_idle & ~ap_sync_kernel_pr_entry98_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                        end
                    end
                    3: begin
                        if (~load_bipedge30_U0.bipedge_stream_blk_n) begin
                            if (~bipedge_stream_0_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_0_V_V_U' written by process 'kernel_pr_kernel_pr.load_value32_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_0_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_0_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_0_V_V_U' read by process 'kernel_pr_kernel_pr.load_value32_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_0_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~load_bipedge30_U0.bipedge_size_out_blk_n) begin
                            if (~bipedge_size_c866_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_size_c866_U' written by process 'kernel_pr_kernel_pr.load_value32_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c866_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_size_c866_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_size_c866_U' read by process 'kernel_pr_kernel_pr.load_value32_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c866_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_bipedge30_U0_ap_ready & load_bipedge30_U0.ap_idle & ~ap_sync_load_value32_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value32_U0'");
                        end
                    end
                    4: begin
                        if (~load_bipedge30_U0.bipedge_stream1_blk_n) begin
                            if (~bipedge_stream_1_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_1_V_V_U' written by process 'kernel_pr_kernel_pr.load_value33_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_1_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_1_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_1_V_V_U' read by process 'kernel_pr_kernel_pr.load_value33_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_1_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~load_bipedge30_U0.bipedge_size_out1_blk_n) begin
                            if (~bipedge_size_c867_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_size_c867_U' written by process 'kernel_pr_kernel_pr.load_value33_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c867_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_size_c867_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_size_c867_U' read by process 'kernel_pr_kernel_pr.load_value33_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c867_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_bipedge30_U0_ap_ready & load_bipedge30_U0.ap_idle & ~ap_sync_load_value33_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value33_U0'");
                        end
                    end
                    5: begin
                        if (~load_bipedge30_U0.bipedge_stream2_blk_n) begin
                            if (~bipedge_stream_2_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_2_V_V_U' written by process 'kernel_pr_kernel_pr.load_value34_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_2_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_2_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_2_V_V_U' read by process 'kernel_pr_kernel_pr.load_value34_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_2_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~load_bipedge30_U0.bipedge_size_out2_blk_n) begin
                            if (~bipedge_size_c868_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_size_c868_U' written by process 'kernel_pr_kernel_pr.load_value34_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c868_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_size_c868_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_size_c868_U' read by process 'kernel_pr_kernel_pr.load_value34_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c868_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_bipedge30_U0_ap_ready & load_bipedge30_U0.ap_idle & ~ap_sync_load_value34_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value34_U0'");
                        end
                    end
                    6: begin
                        if (~load_bipedge30_U0.bipedge_stream3_blk_n) begin
                            if (~bipedge_stream_3_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_3_V_V_U' written by process 'kernel_pr_kernel_pr.load_value35_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_3_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_3_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_3_V_V_U' read by process 'kernel_pr_kernel_pr.load_value35_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_3_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~load_bipedge30_U0.bipedge_size_out3_blk_n) begin
                            if (~bipedge_size_c869_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_size_c869_U' written by process 'kernel_pr_kernel_pr.load_value35_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c869_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_size_c869_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_size_c869_U' read by process 'kernel_pr_kernel_pr.load_value35_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c869_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_bipedge30_U0_ap_ready & load_bipedge30_U0.ap_idle & ~ap_sync_load_value35_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value35_U0'");
                        end
                    end
                    7: begin
                        if (~load_bipedge30_U0.bipedge_stream4_blk_n) begin
                            if (~bipedge_stream_4_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_4_V_V_U' written by process 'kernel_pr_kernel_pr.load_value36_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_4_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_4_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_4_V_V_U' read by process 'kernel_pr_kernel_pr.load_value36_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_4_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~load_bipedge30_U0.bipedge_size_out4_blk_n) begin
                            if (~bipedge_size_c870_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_size_c870_U' written by process 'kernel_pr_kernel_pr.load_value36_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c870_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_size_c870_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_size_c870_U' read by process 'kernel_pr_kernel_pr.load_value36_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c870_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_bipedge30_U0_ap_ready & load_bipedge30_U0.ap_idle & ~ap_sync_load_value36_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value36_U0'");
                        end
                    end
                    8: begin
                        if (~load_bipedge30_U0.bipedge_stream5_blk_n) begin
                            if (~bipedge_stream_5_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_5_V_V_U' written by process 'kernel_pr_kernel_pr.load_value37_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_5_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_5_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_5_V_V_U' read by process 'kernel_pr_kernel_pr.load_value37_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_5_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~load_bipedge30_U0.bipedge_size_out5_blk_n) begin
                            if (~bipedge_size_c871_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_size_c871_U' written by process 'kernel_pr_kernel_pr.load_value37_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c871_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_size_c871_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_size_c871_U' read by process 'kernel_pr_kernel_pr.load_value37_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c871_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_bipedge30_U0_ap_ready & load_bipedge30_U0.ap_idle & ~ap_sync_load_value37_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value37_U0'");
                        end
                    end
                    9: begin
                        if (~load_bipedge30_U0.bipedge_stream6_blk_n) begin
                            if (~bipedge_stream_6_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_6_V_V_U' written by process 'kernel_pr_kernel_pr.load_value38_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_6_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_6_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_6_V_V_U' read by process 'kernel_pr_kernel_pr.load_value38_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_6_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~load_bipedge30_U0.bipedge_size_out6_blk_n) begin
                            if (~bipedge_size_c872_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_size_c872_U' written by process 'kernel_pr_kernel_pr.load_value38_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c872_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_size_c872_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_size_c872_U' read by process 'kernel_pr_kernel_pr.load_value38_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c872_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_bipedge30_U0_ap_ready & load_bipedge30_U0.ap_idle & ~ap_sync_load_value38_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value38_U0'");
                        end
                    end
                    10: begin
                        if (~load_bipedge30_U0.bipedge_stream7_blk_n) begin
                            if (~bipedge_stream_7_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_7_V_V_U' written by process 'kernel_pr_kernel_pr.load_value39_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_7_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_7_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_7_V_V_U' read by process 'kernel_pr_kernel_pr.load_value39_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_7_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~load_bipedge30_U0.bipedge_size_out7_blk_n) begin
                            if (~bipedge_size_c873_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_size_c873_U' written by process 'kernel_pr_kernel_pr.load_value39_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c873_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_size_c873_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_size_c873_U' read by process 'kernel_pr_kernel_pr.load_value39_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c873_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_bipedge30_U0_ap_ready & load_bipedge30_U0.ap_idle & ~ap_sync_load_value39_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value39_U0'");
                        end
                    end
                    2: begin
                        if (ap_sync_load_bipedge30_U0_ap_ready & load_bipedge30_U0.ap_idle & ~ap_sync_load_bipedge31_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge31_U0'");
                        end
                    end
                    11: begin
                        if (ap_sync_load_bipedge30_U0_ap_ready & load_bipedge30_U0.ap_idle & ~ap_sync_load_value40_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value40_U0'");
                        end
                    end
                    12: begin
                        if (ap_sync_load_bipedge30_U0_ap_ready & load_bipedge30_U0.ap_idle & ~ap_sync_load_value41_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value41_U0'");
                        end
                    end
                    13: begin
                        if (ap_sync_load_bipedge30_U0_ap_ready & load_bipedge30_U0.ap_idle & ~ap_sync_load_value42_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value42_U0'");
                        end
                    end
                    14: begin
                        if (ap_sync_load_bipedge30_U0_ap_ready & load_bipedge30_U0.ap_idle & ~ap_sync_load_value43_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value43_U0'");
                        end
                    end
                    15: begin
                        if (ap_sync_load_bipedge30_U0_ap_ready & load_bipedge30_U0.ap_idle & ~ap_sync_load_value44_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value44_U0'");
                        end
                    end
                    16: begin
                        if (ap_sync_load_bipedge30_U0_ap_ready & load_bipedge30_U0.ap_idle & ~ap_sync_load_value45_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value45_U0'");
                        end
                    end
                    17: begin
                        if (ap_sync_load_bipedge30_U0_ap_ready & load_bipedge30_U0.ap_idle & ~ap_sync_load_value46_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value46_U0'");
                        end
                    end
                    18: begin
                        if (ap_sync_load_bipedge30_U0_ap_ready & load_bipedge30_U0.ap_idle & ~ap_sync_load_value47_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value47_U0'");
                        end
                    end
                    endcase
                end
                2 : begin
                    case(index2)
                    0: begin
                        if (~load_bipedge31_U0.bipedge_blk_n) begin
                            if (~hv_bipedge_dram1_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hv_bipedge_dram1_c_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hv_bipedge_dram1_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hv_bipedge_dram1_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hv_bipedge_dram1_c_U' read by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hv_bipedge_dram1_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~load_bipedge31_U0.bipedge_size_blk_n) begin
                            if (~bipedge_size_c865_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_size_c865_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c865_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_size_c865_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_size_c865_U' read by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c865_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_bipedge31_U0_ap_ready & load_bipedge31_U0.ap_idle & ~ap_sync_kernel_pr_entry98_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                        end
                    end
                    11: begin
                        if (~load_bipedge31_U0.bipedge_stream8_blk_n) begin
                            if (~bipedge_stream_8_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_8_V_V_U' written by process 'kernel_pr_kernel_pr.load_value40_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_8_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_8_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_8_V_V_U' read by process 'kernel_pr_kernel_pr.load_value40_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_8_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~load_bipedge31_U0.bipedge_size_out_blk_n) begin
                            if (~bipedge_size_c874_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_size_c874_U' written by process 'kernel_pr_kernel_pr.load_value40_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c874_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_size_c874_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_size_c874_U' read by process 'kernel_pr_kernel_pr.load_value40_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c874_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_bipedge31_U0_ap_ready & load_bipedge31_U0.ap_idle & ~ap_sync_load_value40_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value40_U0'");
                        end
                    end
                    12: begin
                        if (~load_bipedge31_U0.bipedge_stream9_blk_n) begin
                            if (~bipedge_stream_9_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_9_V_V_U' written by process 'kernel_pr_kernel_pr.load_value41_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_9_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_9_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_9_V_V_U' read by process 'kernel_pr_kernel_pr.load_value41_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_9_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~load_bipedge31_U0.bipedge_size_out1_blk_n) begin
                            if (~bipedge_size_c875_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_size_c875_U' written by process 'kernel_pr_kernel_pr.load_value41_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c875_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_size_c875_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_size_c875_U' read by process 'kernel_pr_kernel_pr.load_value41_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c875_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_bipedge31_U0_ap_ready & load_bipedge31_U0.ap_idle & ~ap_sync_load_value41_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value41_U0'");
                        end
                    end
                    13: begin
                        if (~load_bipedge31_U0.bipedge_stream10_blk_n) begin
                            if (~bipedge_stream_10_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_10_V_V_U' written by process 'kernel_pr_kernel_pr.load_value42_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_10_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_10_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_10_V_V_U' read by process 'kernel_pr_kernel_pr.load_value42_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_10_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~load_bipedge31_U0.bipedge_size_out2_blk_n) begin
                            if (~bipedge_size_c876_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_size_c876_U' written by process 'kernel_pr_kernel_pr.load_value42_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c876_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_size_c876_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_size_c876_U' read by process 'kernel_pr_kernel_pr.load_value42_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c876_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_bipedge31_U0_ap_ready & load_bipedge31_U0.ap_idle & ~ap_sync_load_value42_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value42_U0'");
                        end
                    end
                    14: begin
                        if (~load_bipedge31_U0.bipedge_stream11_blk_n) begin
                            if (~bipedge_stream_11_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_11_V_V_U' written by process 'kernel_pr_kernel_pr.load_value43_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_11_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_11_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_11_V_V_U' read by process 'kernel_pr_kernel_pr.load_value43_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_11_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~load_bipedge31_U0.bipedge_size_out3_blk_n) begin
                            if (~bipedge_size_c877_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_size_c877_U' written by process 'kernel_pr_kernel_pr.load_value43_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c877_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_size_c877_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_size_c877_U' read by process 'kernel_pr_kernel_pr.load_value43_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c877_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_bipedge31_U0_ap_ready & load_bipedge31_U0.ap_idle & ~ap_sync_load_value43_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value43_U0'");
                        end
                    end
                    15: begin
                        if (~load_bipedge31_U0.bipedge_stream12_blk_n) begin
                            if (~bipedge_stream_12_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_12_V_V_U' written by process 'kernel_pr_kernel_pr.load_value44_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_12_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_12_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_12_V_V_U' read by process 'kernel_pr_kernel_pr.load_value44_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_12_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~load_bipedge31_U0.bipedge_size_out4_blk_n) begin
                            if (~bipedge_size_c878_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_size_c878_U' written by process 'kernel_pr_kernel_pr.load_value44_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c878_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_size_c878_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_size_c878_U' read by process 'kernel_pr_kernel_pr.load_value44_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c878_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_bipedge31_U0_ap_ready & load_bipedge31_U0.ap_idle & ~ap_sync_load_value44_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value44_U0'");
                        end
                    end
                    16: begin
                        if (~load_bipedge31_U0.bipedge_stream13_blk_n) begin
                            if (~bipedge_stream_13_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_13_V_V_U' written by process 'kernel_pr_kernel_pr.load_value45_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_13_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_13_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_13_V_V_U' read by process 'kernel_pr_kernel_pr.load_value45_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_13_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~load_bipedge31_U0.bipedge_size_out5_blk_n) begin
                            if (~bipedge_size_c879_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_size_c879_U' written by process 'kernel_pr_kernel_pr.load_value45_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c879_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_size_c879_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_size_c879_U' read by process 'kernel_pr_kernel_pr.load_value45_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c879_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_bipedge31_U0_ap_ready & load_bipedge31_U0.ap_idle & ~ap_sync_load_value45_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value45_U0'");
                        end
                    end
                    17: begin
                        if (~load_bipedge31_U0.bipedge_stream14_blk_n) begin
                            if (~bipedge_stream_14_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_14_V_V_U' written by process 'kernel_pr_kernel_pr.load_value46_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_14_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_14_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_14_V_V_U' read by process 'kernel_pr_kernel_pr.load_value46_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_14_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~load_bipedge31_U0.bipedge_size_out6_blk_n) begin
                            if (~bipedge_size_c880_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_size_c880_U' written by process 'kernel_pr_kernel_pr.load_value46_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c880_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_size_c880_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_size_c880_U' read by process 'kernel_pr_kernel_pr.load_value46_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c880_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_bipedge31_U0_ap_ready & load_bipedge31_U0.ap_idle & ~ap_sync_load_value46_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value46_U0'");
                        end
                    end
                    18: begin
                        if (~load_bipedge31_U0.bipedge_stream15_blk_n) begin
                            if (~bipedge_stream_15_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_15_V_V_U' written by process 'kernel_pr_kernel_pr.load_value47_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_15_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_15_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_15_V_V_U' read by process 'kernel_pr_kernel_pr.load_value47_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_15_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~load_bipedge31_U0.bipedge_size_out7_blk_n) begin
                            if (~bipedge_size_c881_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_size_c881_U' written by process 'kernel_pr_kernel_pr.load_value47_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c881_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_size_c881_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_size_c881_U' read by process 'kernel_pr_kernel_pr.load_value47_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c881_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_bipedge31_U0_ap_ready & load_bipedge31_U0.ap_idle & ~ap_sync_load_value47_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value47_U0'");
                        end
                    end
                    1: begin
                        if (ap_sync_load_bipedge31_U0_ap_ready & load_bipedge31_U0.ap_idle & ~ap_sync_load_bipedge30_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge30_U0'");
                        end
                    end
                    3: begin
                        if (ap_sync_load_bipedge31_U0_ap_ready & load_bipedge31_U0.ap_idle & ~ap_sync_load_value32_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value32_U0'");
                        end
                    end
                    4: begin
                        if (ap_sync_load_bipedge31_U0_ap_ready & load_bipedge31_U0.ap_idle & ~ap_sync_load_value33_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value33_U0'");
                        end
                    end
                    5: begin
                        if (ap_sync_load_bipedge31_U0_ap_ready & load_bipedge31_U0.ap_idle & ~ap_sync_load_value34_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value34_U0'");
                        end
                    end
                    6: begin
                        if (ap_sync_load_bipedge31_U0_ap_ready & load_bipedge31_U0.ap_idle & ~ap_sync_load_value35_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value35_U0'");
                        end
                    end
                    7: begin
                        if (ap_sync_load_bipedge31_U0_ap_ready & load_bipedge31_U0.ap_idle & ~ap_sync_load_value36_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value36_U0'");
                        end
                    end
                    8: begin
                        if (ap_sync_load_bipedge31_U0_ap_ready & load_bipedge31_U0.ap_idle & ~ap_sync_load_value37_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value37_U0'");
                        end
                    end
                    9: begin
                        if (ap_sync_load_bipedge31_U0_ap_ready & load_bipedge31_U0.ap_idle & ~ap_sync_load_value38_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value38_U0'");
                        end
                    end
                    10: begin
                        if (ap_sync_load_bipedge31_U0_ap_ready & load_bipedge31_U0.ap_idle & ~ap_sync_load_value39_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value39_U0'");
                        end
                    end
                    endcase
                end
                3 : begin
                    case(index2)
                    0: begin
                        if (~load_value32_U0.value_r_blk_n) begin
                            if (~V_read0_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.V_read0_c_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read0_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~V_read0_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.V_read0_c_U' read by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read0_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_value32_U0_ap_ready & load_value32_U0.ap_idle & ~ap_sync_kernel_pr_entry98_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                        end
                    end
                    1: begin
                        if (~load_value32_U0.bipedge_size_blk_n) begin
                            if (~bipedge_size_c866_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_size_c866_U' written by process 'kernel_pr_kernel_pr.load_bipedge30_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c866_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_size_c866_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_size_c866_U' read by process 'kernel_pr_kernel_pr.load_bipedge30_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c866_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~load_value32_U0.bipedge_stream_V_V_blk_n) begin
                            if (~bipedge_stream_0_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_0_V_V_U' written by process 'kernel_pr_kernel_pr.load_bipedge30_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_0_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_0_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_0_V_V_U' read by process 'kernel_pr_kernel_pr.load_bipedge30_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_0_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_value32_U0_ap_ready & load_value32_U0.ap_idle & ~ap_sync_load_bipedge30_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge30_U0'");
                        end
                    end
                    19: begin
                        if (~load_value32_U0.value_stream_V_V_blk_n) begin
                            if (~value_stream_0_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_0_V_V_U' written by process 'kernel_pr_kernel_pr.write_back48_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_0_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_0_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_0_V_V_U' read by process 'kernel_pr_kernel_pr.write_back48_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_0_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    2: begin
                        if (ap_sync_load_value32_U0_ap_ready & load_value32_U0.ap_idle & ~ap_sync_load_bipedge31_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge31_U0'");
                        end
                    end
                    4: begin
                        if (ap_sync_load_value32_U0_ap_ready & load_value32_U0.ap_idle & ~ap_sync_load_value33_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value33_U0'");
                        end
                    end
                    5: begin
                        if (ap_sync_load_value32_U0_ap_ready & load_value32_U0.ap_idle & ~ap_sync_load_value34_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value34_U0'");
                        end
                    end
                    6: begin
                        if (ap_sync_load_value32_U0_ap_ready & load_value32_U0.ap_idle & ~ap_sync_load_value35_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value35_U0'");
                        end
                    end
                    7: begin
                        if (ap_sync_load_value32_U0_ap_ready & load_value32_U0.ap_idle & ~ap_sync_load_value36_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value36_U0'");
                        end
                    end
                    8: begin
                        if (ap_sync_load_value32_U0_ap_ready & load_value32_U0.ap_idle & ~ap_sync_load_value37_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value37_U0'");
                        end
                    end
                    9: begin
                        if (ap_sync_load_value32_U0_ap_ready & load_value32_U0.ap_idle & ~ap_sync_load_value38_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value38_U0'");
                        end
                    end
                    10: begin
                        if (ap_sync_load_value32_U0_ap_ready & load_value32_U0.ap_idle & ~ap_sync_load_value39_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value39_U0'");
                        end
                    end
                    11: begin
                        if (ap_sync_load_value32_U0_ap_ready & load_value32_U0.ap_idle & ~ap_sync_load_value40_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value40_U0'");
                        end
                    end
                    12: begin
                        if (ap_sync_load_value32_U0_ap_ready & load_value32_U0.ap_idle & ~ap_sync_load_value41_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value41_U0'");
                        end
                    end
                    13: begin
                        if (ap_sync_load_value32_U0_ap_ready & load_value32_U0.ap_idle & ~ap_sync_load_value42_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value42_U0'");
                        end
                    end
                    14: begin
                        if (ap_sync_load_value32_U0_ap_ready & load_value32_U0.ap_idle & ~ap_sync_load_value43_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value43_U0'");
                        end
                    end
                    15: begin
                        if (ap_sync_load_value32_U0_ap_ready & load_value32_U0.ap_idle & ~ap_sync_load_value44_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value44_U0'");
                        end
                    end
                    16: begin
                        if (ap_sync_load_value32_U0_ap_ready & load_value32_U0.ap_idle & ~ap_sync_load_value45_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value45_U0'");
                        end
                    end
                    17: begin
                        if (ap_sync_load_value32_U0_ap_ready & load_value32_U0.ap_idle & ~ap_sync_load_value46_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value46_U0'");
                        end
                    end
                    18: begin
                        if (ap_sync_load_value32_U0_ap_ready & load_value32_U0.ap_idle & ~ap_sync_load_value47_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value47_U0'");
                        end
                    end
                    endcase
                end
                4 : begin
                    case(index2)
                    0: begin
                        if (~load_value33_U0.value_r_blk_n) begin
                            if (~V_read1_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.V_read1_c_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read1_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~V_read1_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.V_read1_c_U' read by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read1_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_value33_U0_ap_ready & load_value33_U0.ap_idle & ~ap_sync_kernel_pr_entry98_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                        end
                    end
                    1: begin
                        if (~load_value33_U0.bipedge_size_blk_n) begin
                            if (~bipedge_size_c867_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_size_c867_U' written by process 'kernel_pr_kernel_pr.load_bipedge30_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c867_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_size_c867_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_size_c867_U' read by process 'kernel_pr_kernel_pr.load_bipedge30_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c867_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~load_value33_U0.bipedge_stream_V_V1_blk_n) begin
                            if (~bipedge_stream_1_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_1_V_V_U' written by process 'kernel_pr_kernel_pr.load_bipedge30_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_1_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_1_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_1_V_V_U' read by process 'kernel_pr_kernel_pr.load_bipedge30_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_1_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_value33_U0_ap_ready & load_value33_U0.ap_idle & ~ap_sync_load_bipedge30_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge30_U0'");
                        end
                    end
                    20: begin
                        if (~load_value33_U0.value_stream_V_V16_blk_n) begin
                            if (~value_stream_1_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_1_V_V_U' written by process 'kernel_pr_kernel_pr.write_back49_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_1_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_1_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_1_V_V_U' read by process 'kernel_pr_kernel_pr.write_back49_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_1_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    2: begin
                        if (ap_sync_load_value33_U0_ap_ready & load_value33_U0.ap_idle & ~ap_sync_load_bipedge31_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge31_U0'");
                        end
                    end
                    3: begin
                        if (ap_sync_load_value33_U0_ap_ready & load_value33_U0.ap_idle & ~ap_sync_load_value32_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value32_U0'");
                        end
                    end
                    5: begin
                        if (ap_sync_load_value33_U0_ap_ready & load_value33_U0.ap_idle & ~ap_sync_load_value34_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value34_U0'");
                        end
                    end
                    6: begin
                        if (ap_sync_load_value33_U0_ap_ready & load_value33_U0.ap_idle & ~ap_sync_load_value35_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value35_U0'");
                        end
                    end
                    7: begin
                        if (ap_sync_load_value33_U0_ap_ready & load_value33_U0.ap_idle & ~ap_sync_load_value36_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value36_U0'");
                        end
                    end
                    8: begin
                        if (ap_sync_load_value33_U0_ap_ready & load_value33_U0.ap_idle & ~ap_sync_load_value37_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value37_U0'");
                        end
                    end
                    9: begin
                        if (ap_sync_load_value33_U0_ap_ready & load_value33_U0.ap_idle & ~ap_sync_load_value38_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value38_U0'");
                        end
                    end
                    10: begin
                        if (ap_sync_load_value33_U0_ap_ready & load_value33_U0.ap_idle & ~ap_sync_load_value39_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value39_U0'");
                        end
                    end
                    11: begin
                        if (ap_sync_load_value33_U0_ap_ready & load_value33_U0.ap_idle & ~ap_sync_load_value40_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value40_U0'");
                        end
                    end
                    12: begin
                        if (ap_sync_load_value33_U0_ap_ready & load_value33_U0.ap_idle & ~ap_sync_load_value41_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value41_U0'");
                        end
                    end
                    13: begin
                        if (ap_sync_load_value33_U0_ap_ready & load_value33_U0.ap_idle & ~ap_sync_load_value42_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value42_U0'");
                        end
                    end
                    14: begin
                        if (ap_sync_load_value33_U0_ap_ready & load_value33_U0.ap_idle & ~ap_sync_load_value43_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value43_U0'");
                        end
                    end
                    15: begin
                        if (ap_sync_load_value33_U0_ap_ready & load_value33_U0.ap_idle & ~ap_sync_load_value44_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value44_U0'");
                        end
                    end
                    16: begin
                        if (ap_sync_load_value33_U0_ap_ready & load_value33_U0.ap_idle & ~ap_sync_load_value45_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value45_U0'");
                        end
                    end
                    17: begin
                        if (ap_sync_load_value33_U0_ap_ready & load_value33_U0.ap_idle & ~ap_sync_load_value46_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value46_U0'");
                        end
                    end
                    18: begin
                        if (ap_sync_load_value33_U0_ap_ready & load_value33_U0.ap_idle & ~ap_sync_load_value47_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value47_U0'");
                        end
                    end
                    endcase
                end
                5 : begin
                    case(index2)
                    0: begin
                        if (~load_value34_U0.value_r_blk_n) begin
                            if (~V_read2_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.V_read2_c_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read2_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~V_read2_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.V_read2_c_U' read by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read2_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_value34_U0_ap_ready & load_value34_U0.ap_idle & ~ap_sync_kernel_pr_entry98_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                        end
                    end
                    1: begin
                        if (~load_value34_U0.bipedge_size_blk_n) begin
                            if (~bipedge_size_c868_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_size_c868_U' written by process 'kernel_pr_kernel_pr.load_bipedge30_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c868_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_size_c868_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_size_c868_U' read by process 'kernel_pr_kernel_pr.load_bipedge30_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c868_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~load_value34_U0.bipedge_stream_V_V2_blk_n) begin
                            if (~bipedge_stream_2_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_2_V_V_U' written by process 'kernel_pr_kernel_pr.load_bipedge30_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_2_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_2_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_2_V_V_U' read by process 'kernel_pr_kernel_pr.load_bipedge30_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_2_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_value34_U0_ap_ready & load_value34_U0.ap_idle & ~ap_sync_load_bipedge30_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge30_U0'");
                        end
                    end
                    21: begin
                        if (~load_value34_U0.value_stream_V_V17_blk_n) begin
                            if (~value_stream_2_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_2_V_V_U' written by process 'kernel_pr_kernel_pr.write_back50_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_2_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_2_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_2_V_V_U' read by process 'kernel_pr_kernel_pr.write_back50_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_2_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    2: begin
                        if (ap_sync_load_value34_U0_ap_ready & load_value34_U0.ap_idle & ~ap_sync_load_bipedge31_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge31_U0'");
                        end
                    end
                    3: begin
                        if (ap_sync_load_value34_U0_ap_ready & load_value34_U0.ap_idle & ~ap_sync_load_value32_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value32_U0'");
                        end
                    end
                    4: begin
                        if (ap_sync_load_value34_U0_ap_ready & load_value34_U0.ap_idle & ~ap_sync_load_value33_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value33_U0'");
                        end
                    end
                    6: begin
                        if (ap_sync_load_value34_U0_ap_ready & load_value34_U0.ap_idle & ~ap_sync_load_value35_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value35_U0'");
                        end
                    end
                    7: begin
                        if (ap_sync_load_value34_U0_ap_ready & load_value34_U0.ap_idle & ~ap_sync_load_value36_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value36_U0'");
                        end
                    end
                    8: begin
                        if (ap_sync_load_value34_U0_ap_ready & load_value34_U0.ap_idle & ~ap_sync_load_value37_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value37_U0'");
                        end
                    end
                    9: begin
                        if (ap_sync_load_value34_U0_ap_ready & load_value34_U0.ap_idle & ~ap_sync_load_value38_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value38_U0'");
                        end
                    end
                    10: begin
                        if (ap_sync_load_value34_U0_ap_ready & load_value34_U0.ap_idle & ~ap_sync_load_value39_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value39_U0'");
                        end
                    end
                    11: begin
                        if (ap_sync_load_value34_U0_ap_ready & load_value34_U0.ap_idle & ~ap_sync_load_value40_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value40_U0'");
                        end
                    end
                    12: begin
                        if (ap_sync_load_value34_U0_ap_ready & load_value34_U0.ap_idle & ~ap_sync_load_value41_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value41_U0'");
                        end
                    end
                    13: begin
                        if (ap_sync_load_value34_U0_ap_ready & load_value34_U0.ap_idle & ~ap_sync_load_value42_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value42_U0'");
                        end
                    end
                    14: begin
                        if (ap_sync_load_value34_U0_ap_ready & load_value34_U0.ap_idle & ~ap_sync_load_value43_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value43_U0'");
                        end
                    end
                    15: begin
                        if (ap_sync_load_value34_U0_ap_ready & load_value34_U0.ap_idle & ~ap_sync_load_value44_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value44_U0'");
                        end
                    end
                    16: begin
                        if (ap_sync_load_value34_U0_ap_ready & load_value34_U0.ap_idle & ~ap_sync_load_value45_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value45_U0'");
                        end
                    end
                    17: begin
                        if (ap_sync_load_value34_U0_ap_ready & load_value34_U0.ap_idle & ~ap_sync_load_value46_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value46_U0'");
                        end
                    end
                    18: begin
                        if (ap_sync_load_value34_U0_ap_ready & load_value34_U0.ap_idle & ~ap_sync_load_value47_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value47_U0'");
                        end
                    end
                    endcase
                end
                6 : begin
                    case(index2)
                    0: begin
                        if (~load_value35_U0.value_r_blk_n) begin
                            if (~V_read3_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.V_read3_c_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read3_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~V_read3_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.V_read3_c_U' read by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read3_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_value35_U0_ap_ready & load_value35_U0.ap_idle & ~ap_sync_kernel_pr_entry98_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                        end
                    end
                    1: begin
                        if (~load_value35_U0.bipedge_size_blk_n) begin
                            if (~bipedge_size_c869_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_size_c869_U' written by process 'kernel_pr_kernel_pr.load_bipedge30_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c869_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_size_c869_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_size_c869_U' read by process 'kernel_pr_kernel_pr.load_bipedge30_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c869_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~load_value35_U0.bipedge_stream_V_V3_blk_n) begin
                            if (~bipedge_stream_3_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_3_V_V_U' written by process 'kernel_pr_kernel_pr.load_bipedge30_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_3_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_3_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_3_V_V_U' read by process 'kernel_pr_kernel_pr.load_bipedge30_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_3_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_value35_U0_ap_ready & load_value35_U0.ap_idle & ~ap_sync_load_bipedge30_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge30_U0'");
                        end
                    end
                    22: begin
                        if (~load_value35_U0.value_stream_V_V18_blk_n) begin
                            if (~value_stream_3_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_3_V_V_U' written by process 'kernel_pr_kernel_pr.write_back51_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_3_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_3_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_3_V_V_U' read by process 'kernel_pr_kernel_pr.write_back51_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_3_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    2: begin
                        if (ap_sync_load_value35_U0_ap_ready & load_value35_U0.ap_idle & ~ap_sync_load_bipedge31_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge31_U0'");
                        end
                    end
                    3: begin
                        if (ap_sync_load_value35_U0_ap_ready & load_value35_U0.ap_idle & ~ap_sync_load_value32_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value32_U0'");
                        end
                    end
                    4: begin
                        if (ap_sync_load_value35_U0_ap_ready & load_value35_U0.ap_idle & ~ap_sync_load_value33_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value33_U0'");
                        end
                    end
                    5: begin
                        if (ap_sync_load_value35_U0_ap_ready & load_value35_U0.ap_idle & ~ap_sync_load_value34_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value34_U0'");
                        end
                    end
                    7: begin
                        if (ap_sync_load_value35_U0_ap_ready & load_value35_U0.ap_idle & ~ap_sync_load_value36_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value36_U0'");
                        end
                    end
                    8: begin
                        if (ap_sync_load_value35_U0_ap_ready & load_value35_U0.ap_idle & ~ap_sync_load_value37_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value37_U0'");
                        end
                    end
                    9: begin
                        if (ap_sync_load_value35_U0_ap_ready & load_value35_U0.ap_idle & ~ap_sync_load_value38_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value38_U0'");
                        end
                    end
                    10: begin
                        if (ap_sync_load_value35_U0_ap_ready & load_value35_U0.ap_idle & ~ap_sync_load_value39_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value39_U0'");
                        end
                    end
                    11: begin
                        if (ap_sync_load_value35_U0_ap_ready & load_value35_U0.ap_idle & ~ap_sync_load_value40_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value40_U0'");
                        end
                    end
                    12: begin
                        if (ap_sync_load_value35_U0_ap_ready & load_value35_U0.ap_idle & ~ap_sync_load_value41_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value41_U0'");
                        end
                    end
                    13: begin
                        if (ap_sync_load_value35_U0_ap_ready & load_value35_U0.ap_idle & ~ap_sync_load_value42_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value42_U0'");
                        end
                    end
                    14: begin
                        if (ap_sync_load_value35_U0_ap_ready & load_value35_U0.ap_idle & ~ap_sync_load_value43_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value43_U0'");
                        end
                    end
                    15: begin
                        if (ap_sync_load_value35_U0_ap_ready & load_value35_U0.ap_idle & ~ap_sync_load_value44_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value44_U0'");
                        end
                    end
                    16: begin
                        if (ap_sync_load_value35_U0_ap_ready & load_value35_U0.ap_idle & ~ap_sync_load_value45_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value45_U0'");
                        end
                    end
                    17: begin
                        if (ap_sync_load_value35_U0_ap_ready & load_value35_U0.ap_idle & ~ap_sync_load_value46_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value46_U0'");
                        end
                    end
                    18: begin
                        if (ap_sync_load_value35_U0_ap_ready & load_value35_U0.ap_idle & ~ap_sync_load_value47_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value47_U0'");
                        end
                    end
                    endcase
                end
                7 : begin
                    case(index2)
                    0: begin
                        if (~load_value36_U0.value_r_blk_n) begin
                            if (~V_read4_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.V_read4_c_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read4_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~V_read4_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.V_read4_c_U' read by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read4_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_value36_U0_ap_ready & load_value36_U0.ap_idle & ~ap_sync_kernel_pr_entry98_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                        end
                    end
                    1: begin
                        if (~load_value36_U0.bipedge_size_blk_n) begin
                            if (~bipedge_size_c870_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_size_c870_U' written by process 'kernel_pr_kernel_pr.load_bipedge30_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c870_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_size_c870_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_size_c870_U' read by process 'kernel_pr_kernel_pr.load_bipedge30_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c870_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~load_value36_U0.bipedge_stream_V_V4_blk_n) begin
                            if (~bipedge_stream_4_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_4_V_V_U' written by process 'kernel_pr_kernel_pr.load_bipedge30_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_4_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_4_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_4_V_V_U' read by process 'kernel_pr_kernel_pr.load_bipedge30_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_4_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_value36_U0_ap_ready & load_value36_U0.ap_idle & ~ap_sync_load_bipedge30_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge30_U0'");
                        end
                    end
                    23: begin
                        if (~load_value36_U0.value_stream_V_V19_blk_n) begin
                            if (~value_stream_4_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_4_V_V_U' written by process 'kernel_pr_kernel_pr.write_back52_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_4_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_4_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_4_V_V_U' read by process 'kernel_pr_kernel_pr.write_back52_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_4_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    2: begin
                        if (ap_sync_load_value36_U0_ap_ready & load_value36_U0.ap_idle & ~ap_sync_load_bipedge31_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge31_U0'");
                        end
                    end
                    3: begin
                        if (ap_sync_load_value36_U0_ap_ready & load_value36_U0.ap_idle & ~ap_sync_load_value32_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value32_U0'");
                        end
                    end
                    4: begin
                        if (ap_sync_load_value36_U0_ap_ready & load_value36_U0.ap_idle & ~ap_sync_load_value33_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value33_U0'");
                        end
                    end
                    5: begin
                        if (ap_sync_load_value36_U0_ap_ready & load_value36_U0.ap_idle & ~ap_sync_load_value34_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value34_U0'");
                        end
                    end
                    6: begin
                        if (ap_sync_load_value36_U0_ap_ready & load_value36_U0.ap_idle & ~ap_sync_load_value35_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value35_U0'");
                        end
                    end
                    8: begin
                        if (ap_sync_load_value36_U0_ap_ready & load_value36_U0.ap_idle & ~ap_sync_load_value37_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value37_U0'");
                        end
                    end
                    9: begin
                        if (ap_sync_load_value36_U0_ap_ready & load_value36_U0.ap_idle & ~ap_sync_load_value38_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value38_U0'");
                        end
                    end
                    10: begin
                        if (ap_sync_load_value36_U0_ap_ready & load_value36_U0.ap_idle & ~ap_sync_load_value39_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value39_U0'");
                        end
                    end
                    11: begin
                        if (ap_sync_load_value36_U0_ap_ready & load_value36_U0.ap_idle & ~ap_sync_load_value40_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value40_U0'");
                        end
                    end
                    12: begin
                        if (ap_sync_load_value36_U0_ap_ready & load_value36_U0.ap_idle & ~ap_sync_load_value41_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value41_U0'");
                        end
                    end
                    13: begin
                        if (ap_sync_load_value36_U0_ap_ready & load_value36_U0.ap_idle & ~ap_sync_load_value42_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value42_U0'");
                        end
                    end
                    14: begin
                        if (ap_sync_load_value36_U0_ap_ready & load_value36_U0.ap_idle & ~ap_sync_load_value43_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value43_U0'");
                        end
                    end
                    15: begin
                        if (ap_sync_load_value36_U0_ap_ready & load_value36_U0.ap_idle & ~ap_sync_load_value44_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value44_U0'");
                        end
                    end
                    16: begin
                        if (ap_sync_load_value36_U0_ap_ready & load_value36_U0.ap_idle & ~ap_sync_load_value45_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value45_U0'");
                        end
                    end
                    17: begin
                        if (ap_sync_load_value36_U0_ap_ready & load_value36_U0.ap_idle & ~ap_sync_load_value46_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value46_U0'");
                        end
                    end
                    18: begin
                        if (ap_sync_load_value36_U0_ap_ready & load_value36_U0.ap_idle & ~ap_sync_load_value47_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value47_U0'");
                        end
                    end
                    endcase
                end
                8 : begin
                    case(index2)
                    0: begin
                        if (~load_value37_U0.value_r_blk_n) begin
                            if (~V_read5_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.V_read5_c_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read5_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~V_read5_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.V_read5_c_U' read by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read5_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_value37_U0_ap_ready & load_value37_U0.ap_idle & ~ap_sync_kernel_pr_entry98_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                        end
                    end
                    1: begin
                        if (~load_value37_U0.bipedge_size_blk_n) begin
                            if (~bipedge_size_c871_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_size_c871_U' written by process 'kernel_pr_kernel_pr.load_bipedge30_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c871_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_size_c871_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_size_c871_U' read by process 'kernel_pr_kernel_pr.load_bipedge30_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c871_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~load_value37_U0.bipedge_stream_V_V5_blk_n) begin
                            if (~bipedge_stream_5_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_5_V_V_U' written by process 'kernel_pr_kernel_pr.load_bipedge30_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_5_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_5_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_5_V_V_U' read by process 'kernel_pr_kernel_pr.load_bipedge30_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_5_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_value37_U0_ap_ready & load_value37_U0.ap_idle & ~ap_sync_load_bipedge30_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge30_U0'");
                        end
                    end
                    24: begin
                        if (~load_value37_U0.value_stream_V_V20_blk_n) begin
                            if (~value_stream_5_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_5_V_V_U' written by process 'kernel_pr_kernel_pr.write_back53_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_5_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_5_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_5_V_V_U' read by process 'kernel_pr_kernel_pr.write_back53_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_5_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    2: begin
                        if (ap_sync_load_value37_U0_ap_ready & load_value37_U0.ap_idle & ~ap_sync_load_bipedge31_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge31_U0'");
                        end
                    end
                    3: begin
                        if (ap_sync_load_value37_U0_ap_ready & load_value37_U0.ap_idle & ~ap_sync_load_value32_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value32_U0'");
                        end
                    end
                    4: begin
                        if (ap_sync_load_value37_U0_ap_ready & load_value37_U0.ap_idle & ~ap_sync_load_value33_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value33_U0'");
                        end
                    end
                    5: begin
                        if (ap_sync_load_value37_U0_ap_ready & load_value37_U0.ap_idle & ~ap_sync_load_value34_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value34_U0'");
                        end
                    end
                    6: begin
                        if (ap_sync_load_value37_U0_ap_ready & load_value37_U0.ap_idle & ~ap_sync_load_value35_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value35_U0'");
                        end
                    end
                    7: begin
                        if (ap_sync_load_value37_U0_ap_ready & load_value37_U0.ap_idle & ~ap_sync_load_value36_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value36_U0'");
                        end
                    end
                    9: begin
                        if (ap_sync_load_value37_U0_ap_ready & load_value37_U0.ap_idle & ~ap_sync_load_value38_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value38_U0'");
                        end
                    end
                    10: begin
                        if (ap_sync_load_value37_U0_ap_ready & load_value37_U0.ap_idle & ~ap_sync_load_value39_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value39_U0'");
                        end
                    end
                    11: begin
                        if (ap_sync_load_value37_U0_ap_ready & load_value37_U0.ap_idle & ~ap_sync_load_value40_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value40_U0'");
                        end
                    end
                    12: begin
                        if (ap_sync_load_value37_U0_ap_ready & load_value37_U0.ap_idle & ~ap_sync_load_value41_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value41_U0'");
                        end
                    end
                    13: begin
                        if (ap_sync_load_value37_U0_ap_ready & load_value37_U0.ap_idle & ~ap_sync_load_value42_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value42_U0'");
                        end
                    end
                    14: begin
                        if (ap_sync_load_value37_U0_ap_ready & load_value37_U0.ap_idle & ~ap_sync_load_value43_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value43_U0'");
                        end
                    end
                    15: begin
                        if (ap_sync_load_value37_U0_ap_ready & load_value37_U0.ap_idle & ~ap_sync_load_value44_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value44_U0'");
                        end
                    end
                    16: begin
                        if (ap_sync_load_value37_U0_ap_ready & load_value37_U0.ap_idle & ~ap_sync_load_value45_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value45_U0'");
                        end
                    end
                    17: begin
                        if (ap_sync_load_value37_U0_ap_ready & load_value37_U0.ap_idle & ~ap_sync_load_value46_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value46_U0'");
                        end
                    end
                    18: begin
                        if (ap_sync_load_value37_U0_ap_ready & load_value37_U0.ap_idle & ~ap_sync_load_value47_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value47_U0'");
                        end
                    end
                    endcase
                end
                9 : begin
                    case(index2)
                    0: begin
                        if (~load_value38_U0.value_r_blk_n) begin
                            if (~V_read6_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.V_read6_c_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read6_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~V_read6_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.V_read6_c_U' read by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read6_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_value38_U0_ap_ready & load_value38_U0.ap_idle & ~ap_sync_kernel_pr_entry98_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                        end
                    end
                    1: begin
                        if (~load_value38_U0.bipedge_size_blk_n) begin
                            if (~bipedge_size_c872_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_size_c872_U' written by process 'kernel_pr_kernel_pr.load_bipedge30_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c872_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_size_c872_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_size_c872_U' read by process 'kernel_pr_kernel_pr.load_bipedge30_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c872_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~load_value38_U0.bipedge_stream_V_V6_blk_n) begin
                            if (~bipedge_stream_6_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_6_V_V_U' written by process 'kernel_pr_kernel_pr.load_bipedge30_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_6_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_6_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_6_V_V_U' read by process 'kernel_pr_kernel_pr.load_bipedge30_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_6_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_value38_U0_ap_ready & load_value38_U0.ap_idle & ~ap_sync_load_bipedge30_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge30_U0'");
                        end
                    end
                    25: begin
                        if (~load_value38_U0.value_stream_V_V21_blk_n) begin
                            if (~value_stream_6_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_6_V_V_U' written by process 'kernel_pr_kernel_pr.write_back54_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_6_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_6_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_6_V_V_U' read by process 'kernel_pr_kernel_pr.write_back54_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_6_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    2: begin
                        if (ap_sync_load_value38_U0_ap_ready & load_value38_U0.ap_idle & ~ap_sync_load_bipedge31_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge31_U0'");
                        end
                    end
                    3: begin
                        if (ap_sync_load_value38_U0_ap_ready & load_value38_U0.ap_idle & ~ap_sync_load_value32_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value32_U0'");
                        end
                    end
                    4: begin
                        if (ap_sync_load_value38_U0_ap_ready & load_value38_U0.ap_idle & ~ap_sync_load_value33_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value33_U0'");
                        end
                    end
                    5: begin
                        if (ap_sync_load_value38_U0_ap_ready & load_value38_U0.ap_idle & ~ap_sync_load_value34_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value34_U0'");
                        end
                    end
                    6: begin
                        if (ap_sync_load_value38_U0_ap_ready & load_value38_U0.ap_idle & ~ap_sync_load_value35_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value35_U0'");
                        end
                    end
                    7: begin
                        if (ap_sync_load_value38_U0_ap_ready & load_value38_U0.ap_idle & ~ap_sync_load_value36_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value36_U0'");
                        end
                    end
                    8: begin
                        if (ap_sync_load_value38_U0_ap_ready & load_value38_U0.ap_idle & ~ap_sync_load_value37_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value37_U0'");
                        end
                    end
                    10: begin
                        if (ap_sync_load_value38_U0_ap_ready & load_value38_U0.ap_idle & ~ap_sync_load_value39_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value39_U0'");
                        end
                    end
                    11: begin
                        if (ap_sync_load_value38_U0_ap_ready & load_value38_U0.ap_idle & ~ap_sync_load_value40_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value40_U0'");
                        end
                    end
                    12: begin
                        if (ap_sync_load_value38_U0_ap_ready & load_value38_U0.ap_idle & ~ap_sync_load_value41_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value41_U0'");
                        end
                    end
                    13: begin
                        if (ap_sync_load_value38_U0_ap_ready & load_value38_U0.ap_idle & ~ap_sync_load_value42_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value42_U0'");
                        end
                    end
                    14: begin
                        if (ap_sync_load_value38_U0_ap_ready & load_value38_U0.ap_idle & ~ap_sync_load_value43_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value43_U0'");
                        end
                    end
                    15: begin
                        if (ap_sync_load_value38_U0_ap_ready & load_value38_U0.ap_idle & ~ap_sync_load_value44_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value44_U0'");
                        end
                    end
                    16: begin
                        if (ap_sync_load_value38_U0_ap_ready & load_value38_U0.ap_idle & ~ap_sync_load_value45_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value45_U0'");
                        end
                    end
                    17: begin
                        if (ap_sync_load_value38_U0_ap_ready & load_value38_U0.ap_idle & ~ap_sync_load_value46_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value46_U0'");
                        end
                    end
                    18: begin
                        if (ap_sync_load_value38_U0_ap_ready & load_value38_U0.ap_idle & ~ap_sync_load_value47_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value47_U0'");
                        end
                    end
                    endcase
                end
                10 : begin
                    case(index2)
                    0: begin
                        if (~load_value39_U0.value_r_blk_n) begin
                            if (~V_read7_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.V_read7_c_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read7_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~V_read7_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.V_read7_c_U' read by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read7_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_value39_U0_ap_ready & load_value39_U0.ap_idle & ~ap_sync_kernel_pr_entry98_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                        end
                    end
                    1: begin
                        if (~load_value39_U0.bipedge_size_blk_n) begin
                            if (~bipedge_size_c873_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_size_c873_U' written by process 'kernel_pr_kernel_pr.load_bipedge30_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c873_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_size_c873_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_size_c873_U' read by process 'kernel_pr_kernel_pr.load_bipedge30_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c873_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~load_value39_U0.bipedge_stream_V_V7_blk_n) begin
                            if (~bipedge_stream_7_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_7_V_V_U' written by process 'kernel_pr_kernel_pr.load_bipedge30_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_7_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_7_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_7_V_V_U' read by process 'kernel_pr_kernel_pr.load_bipedge30_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_7_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_value39_U0_ap_ready & load_value39_U0.ap_idle & ~ap_sync_load_bipedge30_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge30_U0'");
                        end
                    end
                    26: begin
                        if (~load_value39_U0.value_stream_V_V22_blk_n) begin
                            if (~value_stream_7_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_7_V_V_U' written by process 'kernel_pr_kernel_pr.write_back55_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_7_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_7_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_7_V_V_U' read by process 'kernel_pr_kernel_pr.write_back55_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_7_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    2: begin
                        if (ap_sync_load_value39_U0_ap_ready & load_value39_U0.ap_idle & ~ap_sync_load_bipedge31_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge31_U0'");
                        end
                    end
                    3: begin
                        if (ap_sync_load_value39_U0_ap_ready & load_value39_U0.ap_idle & ~ap_sync_load_value32_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value32_U0'");
                        end
                    end
                    4: begin
                        if (ap_sync_load_value39_U0_ap_ready & load_value39_U0.ap_idle & ~ap_sync_load_value33_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value33_U0'");
                        end
                    end
                    5: begin
                        if (ap_sync_load_value39_U0_ap_ready & load_value39_U0.ap_idle & ~ap_sync_load_value34_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value34_U0'");
                        end
                    end
                    6: begin
                        if (ap_sync_load_value39_U0_ap_ready & load_value39_U0.ap_idle & ~ap_sync_load_value35_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value35_U0'");
                        end
                    end
                    7: begin
                        if (ap_sync_load_value39_U0_ap_ready & load_value39_U0.ap_idle & ~ap_sync_load_value36_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value36_U0'");
                        end
                    end
                    8: begin
                        if (ap_sync_load_value39_U0_ap_ready & load_value39_U0.ap_idle & ~ap_sync_load_value37_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value37_U0'");
                        end
                    end
                    9: begin
                        if (ap_sync_load_value39_U0_ap_ready & load_value39_U0.ap_idle & ~ap_sync_load_value38_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value38_U0'");
                        end
                    end
                    11: begin
                        if (ap_sync_load_value39_U0_ap_ready & load_value39_U0.ap_idle & ~ap_sync_load_value40_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value40_U0'");
                        end
                    end
                    12: begin
                        if (ap_sync_load_value39_U0_ap_ready & load_value39_U0.ap_idle & ~ap_sync_load_value41_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value41_U0'");
                        end
                    end
                    13: begin
                        if (ap_sync_load_value39_U0_ap_ready & load_value39_U0.ap_idle & ~ap_sync_load_value42_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value42_U0'");
                        end
                    end
                    14: begin
                        if (ap_sync_load_value39_U0_ap_ready & load_value39_U0.ap_idle & ~ap_sync_load_value43_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value43_U0'");
                        end
                    end
                    15: begin
                        if (ap_sync_load_value39_U0_ap_ready & load_value39_U0.ap_idle & ~ap_sync_load_value44_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value44_U0'");
                        end
                    end
                    16: begin
                        if (ap_sync_load_value39_U0_ap_ready & load_value39_U0.ap_idle & ~ap_sync_load_value45_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value45_U0'");
                        end
                    end
                    17: begin
                        if (ap_sync_load_value39_U0_ap_ready & load_value39_U0.ap_idle & ~ap_sync_load_value46_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value46_U0'");
                        end
                    end
                    18: begin
                        if (ap_sync_load_value39_U0_ap_ready & load_value39_U0.ap_idle & ~ap_sync_load_value47_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value47_U0'");
                        end
                    end
                    endcase
                end
                11 : begin
                    case(index2)
                    0: begin
                        if (~load_value40_U0.value_r_blk_n) begin
                            if (~V_read8_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.V_read8_c_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read8_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~V_read8_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.V_read8_c_U' read by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read8_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_value40_U0_ap_ready & load_value40_U0.ap_idle & ~ap_sync_kernel_pr_entry98_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                        end
                    end
                    2: begin
                        if (~load_value40_U0.bipedge_size_blk_n) begin
                            if (~bipedge_size_c874_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_size_c874_U' written by process 'kernel_pr_kernel_pr.load_bipedge31_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c874_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_size_c874_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_size_c874_U' read by process 'kernel_pr_kernel_pr.load_bipedge31_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c874_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~load_value40_U0.bipedge_stream_V_V8_blk_n) begin
                            if (~bipedge_stream_8_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_8_V_V_U' written by process 'kernel_pr_kernel_pr.load_bipedge31_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_8_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_8_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_8_V_V_U' read by process 'kernel_pr_kernel_pr.load_bipedge31_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_8_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_value40_U0_ap_ready & load_value40_U0.ap_idle & ~ap_sync_load_bipedge31_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge31_U0'");
                        end
                    end
                    27: begin
                        if (~load_value40_U0.value_stream_V_V23_blk_n) begin
                            if (~value_stream_8_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_8_V_V_U' written by process 'kernel_pr_kernel_pr.write_back56_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_8_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_8_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_8_V_V_U' read by process 'kernel_pr_kernel_pr.write_back56_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_8_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    1: begin
                        if (ap_sync_load_value40_U0_ap_ready & load_value40_U0.ap_idle & ~ap_sync_load_bipedge30_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge30_U0'");
                        end
                    end
                    3: begin
                        if (ap_sync_load_value40_U0_ap_ready & load_value40_U0.ap_idle & ~ap_sync_load_value32_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value32_U0'");
                        end
                    end
                    4: begin
                        if (ap_sync_load_value40_U0_ap_ready & load_value40_U0.ap_idle & ~ap_sync_load_value33_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value33_U0'");
                        end
                    end
                    5: begin
                        if (ap_sync_load_value40_U0_ap_ready & load_value40_U0.ap_idle & ~ap_sync_load_value34_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value34_U0'");
                        end
                    end
                    6: begin
                        if (ap_sync_load_value40_U0_ap_ready & load_value40_U0.ap_idle & ~ap_sync_load_value35_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value35_U0'");
                        end
                    end
                    7: begin
                        if (ap_sync_load_value40_U0_ap_ready & load_value40_U0.ap_idle & ~ap_sync_load_value36_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value36_U0'");
                        end
                    end
                    8: begin
                        if (ap_sync_load_value40_U0_ap_ready & load_value40_U0.ap_idle & ~ap_sync_load_value37_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value37_U0'");
                        end
                    end
                    9: begin
                        if (ap_sync_load_value40_U0_ap_ready & load_value40_U0.ap_idle & ~ap_sync_load_value38_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value38_U0'");
                        end
                    end
                    10: begin
                        if (ap_sync_load_value40_U0_ap_ready & load_value40_U0.ap_idle & ~ap_sync_load_value39_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value39_U0'");
                        end
                    end
                    12: begin
                        if (ap_sync_load_value40_U0_ap_ready & load_value40_U0.ap_idle & ~ap_sync_load_value41_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value41_U0'");
                        end
                    end
                    13: begin
                        if (ap_sync_load_value40_U0_ap_ready & load_value40_U0.ap_idle & ~ap_sync_load_value42_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value42_U0'");
                        end
                    end
                    14: begin
                        if (ap_sync_load_value40_U0_ap_ready & load_value40_U0.ap_idle & ~ap_sync_load_value43_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value43_U0'");
                        end
                    end
                    15: begin
                        if (ap_sync_load_value40_U0_ap_ready & load_value40_U0.ap_idle & ~ap_sync_load_value44_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value44_U0'");
                        end
                    end
                    16: begin
                        if (ap_sync_load_value40_U0_ap_ready & load_value40_U0.ap_idle & ~ap_sync_load_value45_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value45_U0'");
                        end
                    end
                    17: begin
                        if (ap_sync_load_value40_U0_ap_ready & load_value40_U0.ap_idle & ~ap_sync_load_value46_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value46_U0'");
                        end
                    end
                    18: begin
                        if (ap_sync_load_value40_U0_ap_ready & load_value40_U0.ap_idle & ~ap_sync_load_value47_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value47_U0'");
                        end
                    end
                    endcase
                end
                12 : begin
                    case(index2)
                    0: begin
                        if (~load_value41_U0.value_r_blk_n) begin
                            if (~V_read9_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.V_read9_c_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read9_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~V_read9_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.V_read9_c_U' read by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read9_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_value41_U0_ap_ready & load_value41_U0.ap_idle & ~ap_sync_kernel_pr_entry98_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                        end
                    end
                    2: begin
                        if (~load_value41_U0.bipedge_size_blk_n) begin
                            if (~bipedge_size_c875_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_size_c875_U' written by process 'kernel_pr_kernel_pr.load_bipedge31_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c875_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_size_c875_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_size_c875_U' read by process 'kernel_pr_kernel_pr.load_bipedge31_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c875_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~load_value41_U0.bipedge_stream_V_V9_blk_n) begin
                            if (~bipedge_stream_9_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_9_V_V_U' written by process 'kernel_pr_kernel_pr.load_bipedge31_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_9_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_9_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_9_V_V_U' read by process 'kernel_pr_kernel_pr.load_bipedge31_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_9_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_value41_U0_ap_ready & load_value41_U0.ap_idle & ~ap_sync_load_bipedge31_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge31_U0'");
                        end
                    end
                    28: begin
                        if (~load_value41_U0.value_stream_V_V24_blk_n) begin
                            if (~value_stream_9_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_9_V_V_U' written by process 'kernel_pr_kernel_pr.write_back57_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_9_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_9_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_9_V_V_U' read by process 'kernel_pr_kernel_pr.write_back57_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_9_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    1: begin
                        if (ap_sync_load_value41_U0_ap_ready & load_value41_U0.ap_idle & ~ap_sync_load_bipedge30_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge30_U0'");
                        end
                    end
                    3: begin
                        if (ap_sync_load_value41_U0_ap_ready & load_value41_U0.ap_idle & ~ap_sync_load_value32_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value32_U0'");
                        end
                    end
                    4: begin
                        if (ap_sync_load_value41_U0_ap_ready & load_value41_U0.ap_idle & ~ap_sync_load_value33_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value33_U0'");
                        end
                    end
                    5: begin
                        if (ap_sync_load_value41_U0_ap_ready & load_value41_U0.ap_idle & ~ap_sync_load_value34_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value34_U0'");
                        end
                    end
                    6: begin
                        if (ap_sync_load_value41_U0_ap_ready & load_value41_U0.ap_idle & ~ap_sync_load_value35_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value35_U0'");
                        end
                    end
                    7: begin
                        if (ap_sync_load_value41_U0_ap_ready & load_value41_U0.ap_idle & ~ap_sync_load_value36_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value36_U0'");
                        end
                    end
                    8: begin
                        if (ap_sync_load_value41_U0_ap_ready & load_value41_U0.ap_idle & ~ap_sync_load_value37_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value37_U0'");
                        end
                    end
                    9: begin
                        if (ap_sync_load_value41_U0_ap_ready & load_value41_U0.ap_idle & ~ap_sync_load_value38_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value38_U0'");
                        end
                    end
                    10: begin
                        if (ap_sync_load_value41_U0_ap_ready & load_value41_U0.ap_idle & ~ap_sync_load_value39_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value39_U0'");
                        end
                    end
                    11: begin
                        if (ap_sync_load_value41_U0_ap_ready & load_value41_U0.ap_idle & ~ap_sync_load_value40_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value40_U0'");
                        end
                    end
                    13: begin
                        if (ap_sync_load_value41_U0_ap_ready & load_value41_U0.ap_idle & ~ap_sync_load_value42_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value42_U0'");
                        end
                    end
                    14: begin
                        if (ap_sync_load_value41_U0_ap_ready & load_value41_U0.ap_idle & ~ap_sync_load_value43_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value43_U0'");
                        end
                    end
                    15: begin
                        if (ap_sync_load_value41_U0_ap_ready & load_value41_U0.ap_idle & ~ap_sync_load_value44_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value44_U0'");
                        end
                    end
                    16: begin
                        if (ap_sync_load_value41_U0_ap_ready & load_value41_U0.ap_idle & ~ap_sync_load_value45_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value45_U0'");
                        end
                    end
                    17: begin
                        if (ap_sync_load_value41_U0_ap_ready & load_value41_U0.ap_idle & ~ap_sync_load_value46_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value46_U0'");
                        end
                    end
                    18: begin
                        if (ap_sync_load_value41_U0_ap_ready & load_value41_U0.ap_idle & ~ap_sync_load_value47_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value47_U0'");
                        end
                    end
                    endcase
                end
                13 : begin
                    case(index2)
                    0: begin
                        if (~load_value42_U0.value_r_blk_n) begin
                            if (~V_read10_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.V_read10_c_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read10_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~V_read10_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.V_read10_c_U' read by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read10_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_value42_U0_ap_ready & load_value42_U0.ap_idle & ~ap_sync_kernel_pr_entry98_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                        end
                    end
                    2: begin
                        if (~load_value42_U0.bipedge_size_blk_n) begin
                            if (~bipedge_size_c876_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_size_c876_U' written by process 'kernel_pr_kernel_pr.load_bipedge31_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c876_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_size_c876_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_size_c876_U' read by process 'kernel_pr_kernel_pr.load_bipedge31_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c876_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~load_value42_U0.bipedge_stream_V_V10_blk_n) begin
                            if (~bipedge_stream_10_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_10_V_V_U' written by process 'kernel_pr_kernel_pr.load_bipedge31_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_10_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_10_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_10_V_V_U' read by process 'kernel_pr_kernel_pr.load_bipedge31_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_10_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_value42_U0_ap_ready & load_value42_U0.ap_idle & ~ap_sync_load_bipedge31_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge31_U0'");
                        end
                    end
                    29: begin
                        if (~load_value42_U0.value_stream_V_V25_blk_n) begin
                            if (~value_stream_10_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_10_V_V_U' written by process 'kernel_pr_kernel_pr.write_back58_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_10_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_10_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_10_V_V_U' read by process 'kernel_pr_kernel_pr.write_back58_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_10_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    1: begin
                        if (ap_sync_load_value42_U0_ap_ready & load_value42_U0.ap_idle & ~ap_sync_load_bipedge30_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge30_U0'");
                        end
                    end
                    3: begin
                        if (ap_sync_load_value42_U0_ap_ready & load_value42_U0.ap_idle & ~ap_sync_load_value32_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value32_U0'");
                        end
                    end
                    4: begin
                        if (ap_sync_load_value42_U0_ap_ready & load_value42_U0.ap_idle & ~ap_sync_load_value33_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value33_U0'");
                        end
                    end
                    5: begin
                        if (ap_sync_load_value42_U0_ap_ready & load_value42_U0.ap_idle & ~ap_sync_load_value34_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value34_U0'");
                        end
                    end
                    6: begin
                        if (ap_sync_load_value42_U0_ap_ready & load_value42_U0.ap_idle & ~ap_sync_load_value35_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value35_U0'");
                        end
                    end
                    7: begin
                        if (ap_sync_load_value42_U0_ap_ready & load_value42_U0.ap_idle & ~ap_sync_load_value36_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value36_U0'");
                        end
                    end
                    8: begin
                        if (ap_sync_load_value42_U0_ap_ready & load_value42_U0.ap_idle & ~ap_sync_load_value37_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value37_U0'");
                        end
                    end
                    9: begin
                        if (ap_sync_load_value42_U0_ap_ready & load_value42_U0.ap_idle & ~ap_sync_load_value38_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value38_U0'");
                        end
                    end
                    10: begin
                        if (ap_sync_load_value42_U0_ap_ready & load_value42_U0.ap_idle & ~ap_sync_load_value39_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value39_U0'");
                        end
                    end
                    11: begin
                        if (ap_sync_load_value42_U0_ap_ready & load_value42_U0.ap_idle & ~ap_sync_load_value40_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value40_U0'");
                        end
                    end
                    12: begin
                        if (ap_sync_load_value42_U0_ap_ready & load_value42_U0.ap_idle & ~ap_sync_load_value41_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value41_U0'");
                        end
                    end
                    14: begin
                        if (ap_sync_load_value42_U0_ap_ready & load_value42_U0.ap_idle & ~ap_sync_load_value43_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value43_U0'");
                        end
                    end
                    15: begin
                        if (ap_sync_load_value42_U0_ap_ready & load_value42_U0.ap_idle & ~ap_sync_load_value44_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value44_U0'");
                        end
                    end
                    16: begin
                        if (ap_sync_load_value42_U0_ap_ready & load_value42_U0.ap_idle & ~ap_sync_load_value45_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value45_U0'");
                        end
                    end
                    17: begin
                        if (ap_sync_load_value42_U0_ap_ready & load_value42_U0.ap_idle & ~ap_sync_load_value46_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value46_U0'");
                        end
                    end
                    18: begin
                        if (ap_sync_load_value42_U0_ap_ready & load_value42_U0.ap_idle & ~ap_sync_load_value47_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value47_U0'");
                        end
                    end
                    endcase
                end
                14 : begin
                    case(index2)
                    0: begin
                        if (~load_value43_U0.value_r_blk_n) begin
                            if (~V_read11_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.V_read11_c_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read11_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~V_read11_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.V_read11_c_U' read by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read11_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_value43_U0_ap_ready & load_value43_U0.ap_idle & ~ap_sync_kernel_pr_entry98_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                        end
                    end
                    2: begin
                        if (~load_value43_U0.bipedge_size_blk_n) begin
                            if (~bipedge_size_c877_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_size_c877_U' written by process 'kernel_pr_kernel_pr.load_bipedge31_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c877_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_size_c877_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_size_c877_U' read by process 'kernel_pr_kernel_pr.load_bipedge31_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c877_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~load_value43_U0.bipedge_stream_V_V11_blk_n) begin
                            if (~bipedge_stream_11_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_11_V_V_U' written by process 'kernel_pr_kernel_pr.load_bipedge31_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_11_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_11_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_11_V_V_U' read by process 'kernel_pr_kernel_pr.load_bipedge31_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_11_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_value43_U0_ap_ready & load_value43_U0.ap_idle & ~ap_sync_load_bipedge31_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge31_U0'");
                        end
                    end
                    30: begin
                        if (~load_value43_U0.value_stream_V_V26_blk_n) begin
                            if (~value_stream_11_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_11_V_V_U' written by process 'kernel_pr_kernel_pr.write_back59_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_11_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_11_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_11_V_V_U' read by process 'kernel_pr_kernel_pr.write_back59_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_11_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    1: begin
                        if (ap_sync_load_value43_U0_ap_ready & load_value43_U0.ap_idle & ~ap_sync_load_bipedge30_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge30_U0'");
                        end
                    end
                    3: begin
                        if (ap_sync_load_value43_U0_ap_ready & load_value43_U0.ap_idle & ~ap_sync_load_value32_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value32_U0'");
                        end
                    end
                    4: begin
                        if (ap_sync_load_value43_U0_ap_ready & load_value43_U0.ap_idle & ~ap_sync_load_value33_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value33_U0'");
                        end
                    end
                    5: begin
                        if (ap_sync_load_value43_U0_ap_ready & load_value43_U0.ap_idle & ~ap_sync_load_value34_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value34_U0'");
                        end
                    end
                    6: begin
                        if (ap_sync_load_value43_U0_ap_ready & load_value43_U0.ap_idle & ~ap_sync_load_value35_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value35_U0'");
                        end
                    end
                    7: begin
                        if (ap_sync_load_value43_U0_ap_ready & load_value43_U0.ap_idle & ~ap_sync_load_value36_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value36_U0'");
                        end
                    end
                    8: begin
                        if (ap_sync_load_value43_U0_ap_ready & load_value43_U0.ap_idle & ~ap_sync_load_value37_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value37_U0'");
                        end
                    end
                    9: begin
                        if (ap_sync_load_value43_U0_ap_ready & load_value43_U0.ap_idle & ~ap_sync_load_value38_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value38_U0'");
                        end
                    end
                    10: begin
                        if (ap_sync_load_value43_U0_ap_ready & load_value43_U0.ap_idle & ~ap_sync_load_value39_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value39_U0'");
                        end
                    end
                    11: begin
                        if (ap_sync_load_value43_U0_ap_ready & load_value43_U0.ap_idle & ~ap_sync_load_value40_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value40_U0'");
                        end
                    end
                    12: begin
                        if (ap_sync_load_value43_U0_ap_ready & load_value43_U0.ap_idle & ~ap_sync_load_value41_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value41_U0'");
                        end
                    end
                    13: begin
                        if (ap_sync_load_value43_U0_ap_ready & load_value43_U0.ap_idle & ~ap_sync_load_value42_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value42_U0'");
                        end
                    end
                    15: begin
                        if (ap_sync_load_value43_U0_ap_ready & load_value43_U0.ap_idle & ~ap_sync_load_value44_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value44_U0'");
                        end
                    end
                    16: begin
                        if (ap_sync_load_value43_U0_ap_ready & load_value43_U0.ap_idle & ~ap_sync_load_value45_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value45_U0'");
                        end
                    end
                    17: begin
                        if (ap_sync_load_value43_U0_ap_ready & load_value43_U0.ap_idle & ~ap_sync_load_value46_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value46_U0'");
                        end
                    end
                    18: begin
                        if (ap_sync_load_value43_U0_ap_ready & load_value43_U0.ap_idle & ~ap_sync_load_value47_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value47_U0'");
                        end
                    end
                    endcase
                end
                15 : begin
                    case(index2)
                    0: begin
                        if (~load_value44_U0.value_r_blk_n) begin
                            if (~V_read12_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.V_read12_c_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read12_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~V_read12_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.V_read12_c_U' read by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read12_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_value44_U0_ap_ready & load_value44_U0.ap_idle & ~ap_sync_kernel_pr_entry98_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                        end
                    end
                    2: begin
                        if (~load_value44_U0.bipedge_size_blk_n) begin
                            if (~bipedge_size_c878_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_size_c878_U' written by process 'kernel_pr_kernel_pr.load_bipedge31_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c878_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_size_c878_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_size_c878_U' read by process 'kernel_pr_kernel_pr.load_bipedge31_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c878_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~load_value44_U0.bipedge_stream_V_V12_blk_n) begin
                            if (~bipedge_stream_12_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_12_V_V_U' written by process 'kernel_pr_kernel_pr.load_bipedge31_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_12_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_12_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_12_V_V_U' read by process 'kernel_pr_kernel_pr.load_bipedge31_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_12_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_value44_U0_ap_ready & load_value44_U0.ap_idle & ~ap_sync_load_bipedge31_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge31_U0'");
                        end
                    end
                    31: begin
                        if (~load_value44_U0.value_stream_V_V27_blk_n) begin
                            if (~value_stream_12_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_12_V_V_U' written by process 'kernel_pr_kernel_pr.write_back60_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_12_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_12_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_12_V_V_U' read by process 'kernel_pr_kernel_pr.write_back60_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_12_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    1: begin
                        if (ap_sync_load_value44_U0_ap_ready & load_value44_U0.ap_idle & ~ap_sync_load_bipedge30_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge30_U0'");
                        end
                    end
                    3: begin
                        if (ap_sync_load_value44_U0_ap_ready & load_value44_U0.ap_idle & ~ap_sync_load_value32_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value32_U0'");
                        end
                    end
                    4: begin
                        if (ap_sync_load_value44_U0_ap_ready & load_value44_U0.ap_idle & ~ap_sync_load_value33_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value33_U0'");
                        end
                    end
                    5: begin
                        if (ap_sync_load_value44_U0_ap_ready & load_value44_U0.ap_idle & ~ap_sync_load_value34_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value34_U0'");
                        end
                    end
                    6: begin
                        if (ap_sync_load_value44_U0_ap_ready & load_value44_U0.ap_idle & ~ap_sync_load_value35_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value35_U0'");
                        end
                    end
                    7: begin
                        if (ap_sync_load_value44_U0_ap_ready & load_value44_U0.ap_idle & ~ap_sync_load_value36_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value36_U0'");
                        end
                    end
                    8: begin
                        if (ap_sync_load_value44_U0_ap_ready & load_value44_U0.ap_idle & ~ap_sync_load_value37_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value37_U0'");
                        end
                    end
                    9: begin
                        if (ap_sync_load_value44_U0_ap_ready & load_value44_U0.ap_idle & ~ap_sync_load_value38_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value38_U0'");
                        end
                    end
                    10: begin
                        if (ap_sync_load_value44_U0_ap_ready & load_value44_U0.ap_idle & ~ap_sync_load_value39_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value39_U0'");
                        end
                    end
                    11: begin
                        if (ap_sync_load_value44_U0_ap_ready & load_value44_U0.ap_idle & ~ap_sync_load_value40_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value40_U0'");
                        end
                    end
                    12: begin
                        if (ap_sync_load_value44_U0_ap_ready & load_value44_U0.ap_idle & ~ap_sync_load_value41_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value41_U0'");
                        end
                    end
                    13: begin
                        if (ap_sync_load_value44_U0_ap_ready & load_value44_U0.ap_idle & ~ap_sync_load_value42_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value42_U0'");
                        end
                    end
                    14: begin
                        if (ap_sync_load_value44_U0_ap_ready & load_value44_U0.ap_idle & ~ap_sync_load_value43_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value43_U0'");
                        end
                    end
                    16: begin
                        if (ap_sync_load_value44_U0_ap_ready & load_value44_U0.ap_idle & ~ap_sync_load_value45_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value45_U0'");
                        end
                    end
                    17: begin
                        if (ap_sync_load_value44_U0_ap_ready & load_value44_U0.ap_idle & ~ap_sync_load_value46_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value46_U0'");
                        end
                    end
                    18: begin
                        if (ap_sync_load_value44_U0_ap_ready & load_value44_U0.ap_idle & ~ap_sync_load_value47_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value47_U0'");
                        end
                    end
                    endcase
                end
                16 : begin
                    case(index2)
                    0: begin
                        if (~load_value45_U0.value_r_blk_n) begin
                            if (~V_read13_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.V_read13_c_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read13_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~V_read13_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.V_read13_c_U' read by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read13_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_value45_U0_ap_ready & load_value45_U0.ap_idle & ~ap_sync_kernel_pr_entry98_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                        end
                    end
                    2: begin
                        if (~load_value45_U0.bipedge_size_blk_n) begin
                            if (~bipedge_size_c879_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_size_c879_U' written by process 'kernel_pr_kernel_pr.load_bipedge31_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c879_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_size_c879_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_size_c879_U' read by process 'kernel_pr_kernel_pr.load_bipedge31_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c879_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~load_value45_U0.bipedge_stream_V_V13_blk_n) begin
                            if (~bipedge_stream_13_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_13_V_V_U' written by process 'kernel_pr_kernel_pr.load_bipedge31_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_13_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_13_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_13_V_V_U' read by process 'kernel_pr_kernel_pr.load_bipedge31_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_13_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_value45_U0_ap_ready & load_value45_U0.ap_idle & ~ap_sync_load_bipedge31_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge31_U0'");
                        end
                    end
                    32: begin
                        if (~load_value45_U0.value_stream_V_V28_blk_n) begin
                            if (~value_stream_13_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_13_V_V_U' written by process 'kernel_pr_kernel_pr.write_back61_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_13_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_13_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_13_V_V_U' read by process 'kernel_pr_kernel_pr.write_back61_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_13_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    1: begin
                        if (ap_sync_load_value45_U0_ap_ready & load_value45_U0.ap_idle & ~ap_sync_load_bipedge30_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge30_U0'");
                        end
                    end
                    3: begin
                        if (ap_sync_load_value45_U0_ap_ready & load_value45_U0.ap_idle & ~ap_sync_load_value32_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value32_U0'");
                        end
                    end
                    4: begin
                        if (ap_sync_load_value45_U0_ap_ready & load_value45_U0.ap_idle & ~ap_sync_load_value33_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value33_U0'");
                        end
                    end
                    5: begin
                        if (ap_sync_load_value45_U0_ap_ready & load_value45_U0.ap_idle & ~ap_sync_load_value34_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value34_U0'");
                        end
                    end
                    6: begin
                        if (ap_sync_load_value45_U0_ap_ready & load_value45_U0.ap_idle & ~ap_sync_load_value35_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value35_U0'");
                        end
                    end
                    7: begin
                        if (ap_sync_load_value45_U0_ap_ready & load_value45_U0.ap_idle & ~ap_sync_load_value36_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value36_U0'");
                        end
                    end
                    8: begin
                        if (ap_sync_load_value45_U0_ap_ready & load_value45_U0.ap_idle & ~ap_sync_load_value37_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value37_U0'");
                        end
                    end
                    9: begin
                        if (ap_sync_load_value45_U0_ap_ready & load_value45_U0.ap_idle & ~ap_sync_load_value38_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value38_U0'");
                        end
                    end
                    10: begin
                        if (ap_sync_load_value45_U0_ap_ready & load_value45_U0.ap_idle & ~ap_sync_load_value39_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value39_U0'");
                        end
                    end
                    11: begin
                        if (ap_sync_load_value45_U0_ap_ready & load_value45_U0.ap_idle & ~ap_sync_load_value40_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value40_U0'");
                        end
                    end
                    12: begin
                        if (ap_sync_load_value45_U0_ap_ready & load_value45_U0.ap_idle & ~ap_sync_load_value41_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value41_U0'");
                        end
                    end
                    13: begin
                        if (ap_sync_load_value45_U0_ap_ready & load_value45_U0.ap_idle & ~ap_sync_load_value42_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value42_U0'");
                        end
                    end
                    14: begin
                        if (ap_sync_load_value45_U0_ap_ready & load_value45_U0.ap_idle & ~ap_sync_load_value43_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value43_U0'");
                        end
                    end
                    15: begin
                        if (ap_sync_load_value45_U0_ap_ready & load_value45_U0.ap_idle & ~ap_sync_load_value44_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value44_U0'");
                        end
                    end
                    17: begin
                        if (ap_sync_load_value45_U0_ap_ready & load_value45_U0.ap_idle & ~ap_sync_load_value46_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value46_U0'");
                        end
                    end
                    18: begin
                        if (ap_sync_load_value45_U0_ap_ready & load_value45_U0.ap_idle & ~ap_sync_load_value47_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value47_U0'");
                        end
                    end
                    endcase
                end
                17 : begin
                    case(index2)
                    0: begin
                        if (~load_value46_U0.value_r_blk_n) begin
                            if (~V_read14_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.V_read14_c_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read14_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~V_read14_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.V_read14_c_U' read by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read14_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_value46_U0_ap_ready & load_value46_U0.ap_idle & ~ap_sync_kernel_pr_entry98_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                        end
                    end
                    2: begin
                        if (~load_value46_U0.bipedge_size_blk_n) begin
                            if (~bipedge_size_c880_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_size_c880_U' written by process 'kernel_pr_kernel_pr.load_bipedge31_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c880_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_size_c880_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_size_c880_U' read by process 'kernel_pr_kernel_pr.load_bipedge31_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c880_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~load_value46_U0.bipedge_stream_V_V14_blk_n) begin
                            if (~bipedge_stream_14_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_14_V_V_U' written by process 'kernel_pr_kernel_pr.load_bipedge31_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_14_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_14_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_14_V_V_U' read by process 'kernel_pr_kernel_pr.load_bipedge31_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_14_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_value46_U0_ap_ready & load_value46_U0.ap_idle & ~ap_sync_load_bipedge31_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge31_U0'");
                        end
                    end
                    33: begin
                        if (~load_value46_U0.value_stream_V_V29_blk_n) begin
                            if (~value_stream_14_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_14_V_V_U' written by process 'kernel_pr_kernel_pr.write_back62_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_14_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_14_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_14_V_V_U' read by process 'kernel_pr_kernel_pr.write_back62_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_14_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    1: begin
                        if (ap_sync_load_value46_U0_ap_ready & load_value46_U0.ap_idle & ~ap_sync_load_bipedge30_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge30_U0'");
                        end
                    end
                    3: begin
                        if (ap_sync_load_value46_U0_ap_ready & load_value46_U0.ap_idle & ~ap_sync_load_value32_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value32_U0'");
                        end
                    end
                    4: begin
                        if (ap_sync_load_value46_U0_ap_ready & load_value46_U0.ap_idle & ~ap_sync_load_value33_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value33_U0'");
                        end
                    end
                    5: begin
                        if (ap_sync_load_value46_U0_ap_ready & load_value46_U0.ap_idle & ~ap_sync_load_value34_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value34_U0'");
                        end
                    end
                    6: begin
                        if (ap_sync_load_value46_U0_ap_ready & load_value46_U0.ap_idle & ~ap_sync_load_value35_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value35_U0'");
                        end
                    end
                    7: begin
                        if (ap_sync_load_value46_U0_ap_ready & load_value46_U0.ap_idle & ~ap_sync_load_value36_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value36_U0'");
                        end
                    end
                    8: begin
                        if (ap_sync_load_value46_U0_ap_ready & load_value46_U0.ap_idle & ~ap_sync_load_value37_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value37_U0'");
                        end
                    end
                    9: begin
                        if (ap_sync_load_value46_U0_ap_ready & load_value46_U0.ap_idle & ~ap_sync_load_value38_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value38_U0'");
                        end
                    end
                    10: begin
                        if (ap_sync_load_value46_U0_ap_ready & load_value46_U0.ap_idle & ~ap_sync_load_value39_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value39_U0'");
                        end
                    end
                    11: begin
                        if (ap_sync_load_value46_U0_ap_ready & load_value46_U0.ap_idle & ~ap_sync_load_value40_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value40_U0'");
                        end
                    end
                    12: begin
                        if (ap_sync_load_value46_U0_ap_ready & load_value46_U0.ap_idle & ~ap_sync_load_value41_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value41_U0'");
                        end
                    end
                    13: begin
                        if (ap_sync_load_value46_U0_ap_ready & load_value46_U0.ap_idle & ~ap_sync_load_value42_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value42_U0'");
                        end
                    end
                    14: begin
                        if (ap_sync_load_value46_U0_ap_ready & load_value46_U0.ap_idle & ~ap_sync_load_value43_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value43_U0'");
                        end
                    end
                    15: begin
                        if (ap_sync_load_value46_U0_ap_ready & load_value46_U0.ap_idle & ~ap_sync_load_value44_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value44_U0'");
                        end
                    end
                    16: begin
                        if (ap_sync_load_value46_U0_ap_ready & load_value46_U0.ap_idle & ~ap_sync_load_value45_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value45_U0'");
                        end
                    end
                    18: begin
                        if (ap_sync_load_value46_U0_ap_ready & load_value46_U0.ap_idle & ~ap_sync_load_value47_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value47_U0'");
                        end
                    end
                    endcase
                end
                18 : begin
                    case(index2)
                    0: begin
                        if (~load_value47_U0.value_r_blk_n) begin
                            if (~V_read15_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.V_read15_c_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read15_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~V_read15_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.V_read15_c_U' read by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.V_read15_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_value47_U0_ap_ready & load_value47_U0.ap_idle & ~ap_sync_kernel_pr_entry98_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                        end
                    end
                    2: begin
                        if (~load_value47_U0.bipedge_size_blk_n) begin
                            if (~bipedge_size_c881_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_size_c881_U' written by process 'kernel_pr_kernel_pr.load_bipedge31_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c881_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_size_c881_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_size_c881_U' read by process 'kernel_pr_kernel_pr.load_bipedge31_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_size_c881_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~load_value47_U0.bipedge_stream_V_V15_blk_n) begin
                            if (~bipedge_stream_15_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.bipedge_stream_15_V_V_U' written by process 'kernel_pr_kernel_pr.load_bipedge31_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_15_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~bipedge_stream_15_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.bipedge_stream_15_V_V_U' read by process 'kernel_pr_kernel_pr.load_bipedge31_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.bipedge_stream_15_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (ap_sync_load_value47_U0_ap_ready & load_value47_U0.ap_idle & ~ap_sync_load_bipedge31_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge31_U0'");
                        end
                    end
                    34: begin
                        if (~load_value47_U0.value_stream_V_V30_blk_n) begin
                            if (~value_stream_15_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_15_V_V_U' written by process 'kernel_pr_kernel_pr.write_back63_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_15_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_15_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_15_V_V_U' read by process 'kernel_pr_kernel_pr.write_back63_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_15_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    1: begin
                        if (ap_sync_load_value47_U0_ap_ready & load_value47_U0.ap_idle & ~ap_sync_load_bipedge30_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_bipedge30_U0'");
                        end
                    end
                    3: begin
                        if (ap_sync_load_value47_U0_ap_ready & load_value47_U0.ap_idle & ~ap_sync_load_value32_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value32_U0'");
                        end
                    end
                    4: begin
                        if (ap_sync_load_value47_U0_ap_ready & load_value47_U0.ap_idle & ~ap_sync_load_value33_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value33_U0'");
                        end
                    end
                    5: begin
                        if (ap_sync_load_value47_U0_ap_ready & load_value47_U0.ap_idle & ~ap_sync_load_value34_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value34_U0'");
                        end
                    end
                    6: begin
                        if (ap_sync_load_value47_U0_ap_ready & load_value47_U0.ap_idle & ~ap_sync_load_value35_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value35_U0'");
                        end
                    end
                    7: begin
                        if (ap_sync_load_value47_U0_ap_ready & load_value47_U0.ap_idle & ~ap_sync_load_value36_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value36_U0'");
                        end
                    end
                    8: begin
                        if (ap_sync_load_value47_U0_ap_ready & load_value47_U0.ap_idle & ~ap_sync_load_value37_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value37_U0'");
                        end
                    end
                    9: begin
                        if (ap_sync_load_value47_U0_ap_ready & load_value47_U0.ap_idle & ~ap_sync_load_value38_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value38_U0'");
                        end
                    end
                    10: begin
                        if (ap_sync_load_value47_U0_ap_ready & load_value47_U0.ap_idle & ~ap_sync_load_value39_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value39_U0'");
                        end
                    end
                    11: begin
                        if (ap_sync_load_value47_U0_ap_ready & load_value47_U0.ap_idle & ~ap_sync_load_value40_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value40_U0'");
                        end
                    end
                    12: begin
                        if (ap_sync_load_value47_U0_ap_ready & load_value47_U0.ap_idle & ~ap_sync_load_value41_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value41_U0'");
                        end
                    end
                    13: begin
                        if (ap_sync_load_value47_U0_ap_ready & load_value47_U0.ap_idle & ~ap_sync_load_value42_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value42_U0'");
                        end
                    end
                    14: begin
                        if (ap_sync_load_value47_U0_ap_ready & load_value47_U0.ap_idle & ~ap_sync_load_value43_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value43_U0'");
                        end
                    end
                    15: begin
                        if (ap_sync_load_value47_U0_ap_ready & load_value47_U0.ap_idle & ~ap_sync_load_value44_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value44_U0'");
                        end
                    end
                    16: begin
                        if (ap_sync_load_value47_U0_ap_ready & load_value47_U0.ap_idle & ~ap_sync_load_value45_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value45_U0'");
                        end
                    end
                    17: begin
                        if (ap_sync_load_value47_U0_ap_ready & load_value47_U0.ap_idle & ~ap_sync_load_value46_U0_ap_ready) begin
                            $display("//      Blocked by input sync logic with process : 'kernel_pr_kernel_pr.load_value46_U0'");
                        end
                    end
                    endcase
                end
                19 : begin
                    case(index2)
                    0: begin
                        if (~write_back48_U0.H_blk_n) begin
                            if (~H_write0_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write0_c_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write0_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write0_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write0_c_U' read by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write0_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~write_back48_U0.hyperedge_size_blk_n) begin
                            if (~hyperedge_size_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c_U' read by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back48_U0_U.if_empty_n & write_back48_U0.ap_idle & ~start_for_write_back48_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back48_U0_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0',");
                        end
                    end
                    3: begin
                        if (~write_back48_U0.value_stream_V_V_blk_n) begin
                            if (~value_stream_0_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_0_V_V_U' written by process 'kernel_pr_kernel_pr.load_value32_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_0_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_0_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_0_V_V_U' read by process 'kernel_pr_kernel_pr.load_value32_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_0_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    20: begin
                        if (ap_done_reg_0 & write_back48_U0.ap_done & ~write_back49_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back49_U0'");
                        end
                    end
                    21: begin
                        if (ap_done_reg_0 & write_back48_U0.ap_done & ~write_back50_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back50_U0'");
                        end
                    end
                    22: begin
                        if (ap_done_reg_0 & write_back48_U0.ap_done & ~write_back51_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back51_U0'");
                        end
                    end
                    23: begin
                        if (ap_done_reg_0 & write_back48_U0.ap_done & ~write_back52_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back52_U0'");
                        end
                    end
                    24: begin
                        if (ap_done_reg_0 & write_back48_U0.ap_done & ~write_back53_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back53_U0'");
                        end
                    end
                    25: begin
                        if (ap_done_reg_0 & write_back48_U0.ap_done & ~write_back54_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back54_U0'");
                        end
                    end
                    26: begin
                        if (ap_done_reg_0 & write_back48_U0.ap_done & ~write_back55_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back55_U0'");
                        end
                    end
                    27: begin
                        if (ap_done_reg_0 & write_back48_U0.ap_done & ~write_back56_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back56_U0'");
                        end
                    end
                    28: begin
                        if (ap_done_reg_0 & write_back48_U0.ap_done & ~write_back57_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back57_U0'");
                        end
                    end
                    29: begin
                        if (ap_done_reg_0 & write_back48_U0.ap_done & ~write_back58_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back58_U0'");
                        end
                    end
                    30: begin
                        if (ap_done_reg_0 & write_back48_U0.ap_done & ~write_back59_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back59_U0'");
                        end
                    end
                    31: begin
                        if (ap_done_reg_0 & write_back48_U0.ap_done & ~write_back60_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back60_U0'");
                        end
                    end
                    32: begin
                        if (ap_done_reg_0 & write_back48_U0.ap_done & ~write_back61_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back61_U0'");
                        end
                    end
                    33: begin
                        if (ap_done_reg_0 & write_back48_U0.ap_done & ~write_back62_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back62_U0'");
                        end
                    end
                    34: begin
                        if (ap_done_reg_0 & write_back48_U0.ap_done & ~write_back63_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back63_U0'");
                        end
                    end
                    endcase
                end
                20 : begin
                    case(index2)
                    0: begin
                        if (~write_back49_U0.H_blk_n) begin
                            if (~H_write1_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write1_c_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write1_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write1_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write1_c_U' read by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write1_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~write_back49_U0.hyperedge_size_blk_n) begin
                            if (~hyperedge_size_c850_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c850_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c850_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c850_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c850_U' read by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c850_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back49_U0_U.if_empty_n & write_back49_U0.ap_idle & ~start_for_write_back49_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back49_U0_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0',");
                        end
                    end
                    4: begin
                        if (~write_back49_U0.value_stream_V_V1_blk_n) begin
                            if (~value_stream_1_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_1_V_V_U' written by process 'kernel_pr_kernel_pr.load_value33_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_1_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_1_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_1_V_V_U' read by process 'kernel_pr_kernel_pr.load_value33_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_1_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    19: begin
                        if (ap_done_reg_1 & write_back49_U0.ap_done & ~write_back48_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back48_U0'");
                        end
                    end
                    21: begin
                        if (ap_done_reg_1 & write_back49_U0.ap_done & ~write_back50_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back50_U0'");
                        end
                    end
                    22: begin
                        if (ap_done_reg_1 & write_back49_U0.ap_done & ~write_back51_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back51_U0'");
                        end
                    end
                    23: begin
                        if (ap_done_reg_1 & write_back49_U0.ap_done & ~write_back52_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back52_U0'");
                        end
                    end
                    24: begin
                        if (ap_done_reg_1 & write_back49_U0.ap_done & ~write_back53_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back53_U0'");
                        end
                    end
                    25: begin
                        if (ap_done_reg_1 & write_back49_U0.ap_done & ~write_back54_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back54_U0'");
                        end
                    end
                    26: begin
                        if (ap_done_reg_1 & write_back49_U0.ap_done & ~write_back55_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back55_U0'");
                        end
                    end
                    27: begin
                        if (ap_done_reg_1 & write_back49_U0.ap_done & ~write_back56_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back56_U0'");
                        end
                    end
                    28: begin
                        if (ap_done_reg_1 & write_back49_U0.ap_done & ~write_back57_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back57_U0'");
                        end
                    end
                    29: begin
                        if (ap_done_reg_1 & write_back49_U0.ap_done & ~write_back58_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back58_U0'");
                        end
                    end
                    30: begin
                        if (ap_done_reg_1 & write_back49_U0.ap_done & ~write_back59_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back59_U0'");
                        end
                    end
                    31: begin
                        if (ap_done_reg_1 & write_back49_U0.ap_done & ~write_back60_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back60_U0'");
                        end
                    end
                    32: begin
                        if (ap_done_reg_1 & write_back49_U0.ap_done & ~write_back61_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back61_U0'");
                        end
                    end
                    33: begin
                        if (ap_done_reg_1 & write_back49_U0.ap_done & ~write_back62_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back62_U0'");
                        end
                    end
                    34: begin
                        if (ap_done_reg_1 & write_back49_U0.ap_done & ~write_back63_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back63_U0'");
                        end
                    end
                    endcase
                end
                21 : begin
                    case(index2)
                    0: begin
                        if (~write_back50_U0.H_blk_n) begin
                            if (~H_write2_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write2_c_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write2_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write2_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write2_c_U' read by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write2_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~write_back50_U0.hyperedge_size_blk_n) begin
                            if (~hyperedge_size_c851_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c851_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c851_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c851_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c851_U' read by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c851_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back50_U0_U.if_empty_n & write_back50_U0.ap_idle & ~start_for_write_back50_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back50_U0_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0',");
                        end
                    end
                    5: begin
                        if (~write_back50_U0.value_stream_V_V2_blk_n) begin
                            if (~value_stream_2_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_2_V_V_U' written by process 'kernel_pr_kernel_pr.load_value34_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_2_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_2_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_2_V_V_U' read by process 'kernel_pr_kernel_pr.load_value34_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_2_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    19: begin
                        if (ap_done_reg_2 & write_back50_U0.ap_done & ~write_back48_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back48_U0'");
                        end
                    end
                    20: begin
                        if (ap_done_reg_2 & write_back50_U0.ap_done & ~write_back49_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back49_U0'");
                        end
                    end
                    22: begin
                        if (ap_done_reg_2 & write_back50_U0.ap_done & ~write_back51_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back51_U0'");
                        end
                    end
                    23: begin
                        if (ap_done_reg_2 & write_back50_U0.ap_done & ~write_back52_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back52_U0'");
                        end
                    end
                    24: begin
                        if (ap_done_reg_2 & write_back50_U0.ap_done & ~write_back53_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back53_U0'");
                        end
                    end
                    25: begin
                        if (ap_done_reg_2 & write_back50_U0.ap_done & ~write_back54_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back54_U0'");
                        end
                    end
                    26: begin
                        if (ap_done_reg_2 & write_back50_U0.ap_done & ~write_back55_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back55_U0'");
                        end
                    end
                    27: begin
                        if (ap_done_reg_2 & write_back50_U0.ap_done & ~write_back56_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back56_U0'");
                        end
                    end
                    28: begin
                        if (ap_done_reg_2 & write_back50_U0.ap_done & ~write_back57_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back57_U0'");
                        end
                    end
                    29: begin
                        if (ap_done_reg_2 & write_back50_U0.ap_done & ~write_back58_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back58_U0'");
                        end
                    end
                    30: begin
                        if (ap_done_reg_2 & write_back50_U0.ap_done & ~write_back59_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back59_U0'");
                        end
                    end
                    31: begin
                        if (ap_done_reg_2 & write_back50_U0.ap_done & ~write_back60_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back60_U0'");
                        end
                    end
                    32: begin
                        if (ap_done_reg_2 & write_back50_U0.ap_done & ~write_back61_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back61_U0'");
                        end
                    end
                    33: begin
                        if (ap_done_reg_2 & write_back50_U0.ap_done & ~write_back62_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back62_U0'");
                        end
                    end
                    34: begin
                        if (ap_done_reg_2 & write_back50_U0.ap_done & ~write_back63_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back63_U0'");
                        end
                    end
                    endcase
                end
                22 : begin
                    case(index2)
                    0: begin
                        if (~write_back51_U0.H_blk_n) begin
                            if (~H_write3_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write3_c_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write3_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write3_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write3_c_U' read by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write3_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~write_back51_U0.hyperedge_size_blk_n) begin
                            if (~hyperedge_size_c852_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c852_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c852_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c852_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c852_U' read by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c852_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back51_U0_U.if_empty_n & write_back51_U0.ap_idle & ~start_for_write_back51_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back51_U0_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0',");
                        end
                    end
                    6: begin
                        if (~write_back51_U0.value_stream_V_V3_blk_n) begin
                            if (~value_stream_3_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_3_V_V_U' written by process 'kernel_pr_kernel_pr.load_value35_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_3_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_3_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_3_V_V_U' read by process 'kernel_pr_kernel_pr.load_value35_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_3_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    19: begin
                        if (ap_done_reg_3 & write_back51_U0.ap_done & ~write_back48_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back48_U0'");
                        end
                    end
                    20: begin
                        if (ap_done_reg_3 & write_back51_U0.ap_done & ~write_back49_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back49_U0'");
                        end
                    end
                    21: begin
                        if (ap_done_reg_3 & write_back51_U0.ap_done & ~write_back50_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back50_U0'");
                        end
                    end
                    23: begin
                        if (ap_done_reg_3 & write_back51_U0.ap_done & ~write_back52_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back52_U0'");
                        end
                    end
                    24: begin
                        if (ap_done_reg_3 & write_back51_U0.ap_done & ~write_back53_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back53_U0'");
                        end
                    end
                    25: begin
                        if (ap_done_reg_3 & write_back51_U0.ap_done & ~write_back54_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back54_U0'");
                        end
                    end
                    26: begin
                        if (ap_done_reg_3 & write_back51_U0.ap_done & ~write_back55_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back55_U0'");
                        end
                    end
                    27: begin
                        if (ap_done_reg_3 & write_back51_U0.ap_done & ~write_back56_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back56_U0'");
                        end
                    end
                    28: begin
                        if (ap_done_reg_3 & write_back51_U0.ap_done & ~write_back57_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back57_U0'");
                        end
                    end
                    29: begin
                        if (ap_done_reg_3 & write_back51_U0.ap_done & ~write_back58_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back58_U0'");
                        end
                    end
                    30: begin
                        if (ap_done_reg_3 & write_back51_U0.ap_done & ~write_back59_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back59_U0'");
                        end
                    end
                    31: begin
                        if (ap_done_reg_3 & write_back51_U0.ap_done & ~write_back60_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back60_U0'");
                        end
                    end
                    32: begin
                        if (ap_done_reg_3 & write_back51_U0.ap_done & ~write_back61_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back61_U0'");
                        end
                    end
                    33: begin
                        if (ap_done_reg_3 & write_back51_U0.ap_done & ~write_back62_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back62_U0'");
                        end
                    end
                    34: begin
                        if (ap_done_reg_3 & write_back51_U0.ap_done & ~write_back63_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back63_U0'");
                        end
                    end
                    endcase
                end
                23 : begin
                    case(index2)
                    0: begin
                        if (~write_back52_U0.H_blk_n) begin
                            if (~H_write4_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write4_c_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write4_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write4_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write4_c_U' read by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write4_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~write_back52_U0.hyperedge_size_blk_n) begin
                            if (~hyperedge_size_c853_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c853_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c853_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c853_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c853_U' read by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c853_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back52_U0_U.if_empty_n & write_back52_U0.ap_idle & ~start_for_write_back52_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back52_U0_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0',");
                        end
                    end
                    7: begin
                        if (~write_back52_U0.value_stream_V_V4_blk_n) begin
                            if (~value_stream_4_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_4_V_V_U' written by process 'kernel_pr_kernel_pr.load_value36_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_4_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_4_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_4_V_V_U' read by process 'kernel_pr_kernel_pr.load_value36_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_4_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    19: begin
                        if (ap_done_reg_4 & write_back52_U0.ap_done & ~write_back48_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back48_U0'");
                        end
                    end
                    20: begin
                        if (ap_done_reg_4 & write_back52_U0.ap_done & ~write_back49_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back49_U0'");
                        end
                    end
                    21: begin
                        if (ap_done_reg_4 & write_back52_U0.ap_done & ~write_back50_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back50_U0'");
                        end
                    end
                    22: begin
                        if (ap_done_reg_4 & write_back52_U0.ap_done & ~write_back51_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back51_U0'");
                        end
                    end
                    24: begin
                        if (ap_done_reg_4 & write_back52_U0.ap_done & ~write_back53_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back53_U0'");
                        end
                    end
                    25: begin
                        if (ap_done_reg_4 & write_back52_U0.ap_done & ~write_back54_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back54_U0'");
                        end
                    end
                    26: begin
                        if (ap_done_reg_4 & write_back52_U0.ap_done & ~write_back55_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back55_U0'");
                        end
                    end
                    27: begin
                        if (ap_done_reg_4 & write_back52_U0.ap_done & ~write_back56_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back56_U0'");
                        end
                    end
                    28: begin
                        if (ap_done_reg_4 & write_back52_U0.ap_done & ~write_back57_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back57_U0'");
                        end
                    end
                    29: begin
                        if (ap_done_reg_4 & write_back52_U0.ap_done & ~write_back58_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back58_U0'");
                        end
                    end
                    30: begin
                        if (ap_done_reg_4 & write_back52_U0.ap_done & ~write_back59_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back59_U0'");
                        end
                    end
                    31: begin
                        if (ap_done_reg_4 & write_back52_U0.ap_done & ~write_back60_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back60_U0'");
                        end
                    end
                    32: begin
                        if (ap_done_reg_4 & write_back52_U0.ap_done & ~write_back61_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back61_U0'");
                        end
                    end
                    33: begin
                        if (ap_done_reg_4 & write_back52_U0.ap_done & ~write_back62_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back62_U0'");
                        end
                    end
                    34: begin
                        if (ap_done_reg_4 & write_back52_U0.ap_done & ~write_back63_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back63_U0'");
                        end
                    end
                    endcase
                end
                24 : begin
                    case(index2)
                    0: begin
                        if (~write_back53_U0.H_blk_n) begin
                            if (~H_write5_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write5_c_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write5_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write5_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write5_c_U' read by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write5_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~write_back53_U0.hyperedge_size_blk_n) begin
                            if (~hyperedge_size_c854_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c854_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c854_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c854_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c854_U' read by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c854_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back53_U0_U.if_empty_n & write_back53_U0.ap_idle & ~start_for_write_back53_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back53_U0_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0',");
                        end
                    end
                    8: begin
                        if (~write_back53_U0.value_stream_V_V5_blk_n) begin
                            if (~value_stream_5_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_5_V_V_U' written by process 'kernel_pr_kernel_pr.load_value37_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_5_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_5_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_5_V_V_U' read by process 'kernel_pr_kernel_pr.load_value37_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_5_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    19: begin
                        if (ap_done_reg_5 & write_back53_U0.ap_done & ~write_back48_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back48_U0'");
                        end
                    end
                    20: begin
                        if (ap_done_reg_5 & write_back53_U0.ap_done & ~write_back49_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back49_U0'");
                        end
                    end
                    21: begin
                        if (ap_done_reg_5 & write_back53_U0.ap_done & ~write_back50_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back50_U0'");
                        end
                    end
                    22: begin
                        if (ap_done_reg_5 & write_back53_U0.ap_done & ~write_back51_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back51_U0'");
                        end
                    end
                    23: begin
                        if (ap_done_reg_5 & write_back53_U0.ap_done & ~write_back52_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back52_U0'");
                        end
                    end
                    25: begin
                        if (ap_done_reg_5 & write_back53_U0.ap_done & ~write_back54_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back54_U0'");
                        end
                    end
                    26: begin
                        if (ap_done_reg_5 & write_back53_U0.ap_done & ~write_back55_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back55_U0'");
                        end
                    end
                    27: begin
                        if (ap_done_reg_5 & write_back53_U0.ap_done & ~write_back56_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back56_U0'");
                        end
                    end
                    28: begin
                        if (ap_done_reg_5 & write_back53_U0.ap_done & ~write_back57_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back57_U0'");
                        end
                    end
                    29: begin
                        if (ap_done_reg_5 & write_back53_U0.ap_done & ~write_back58_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back58_U0'");
                        end
                    end
                    30: begin
                        if (ap_done_reg_5 & write_back53_U0.ap_done & ~write_back59_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back59_U0'");
                        end
                    end
                    31: begin
                        if (ap_done_reg_5 & write_back53_U0.ap_done & ~write_back60_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back60_U0'");
                        end
                    end
                    32: begin
                        if (ap_done_reg_5 & write_back53_U0.ap_done & ~write_back61_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back61_U0'");
                        end
                    end
                    33: begin
                        if (ap_done_reg_5 & write_back53_U0.ap_done & ~write_back62_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back62_U0'");
                        end
                    end
                    34: begin
                        if (ap_done_reg_5 & write_back53_U0.ap_done & ~write_back63_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back63_U0'");
                        end
                    end
                    endcase
                end
                25 : begin
                    case(index2)
                    0: begin
                        if (~write_back54_U0.H_blk_n) begin
                            if (~H_write6_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write6_c_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write6_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write6_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write6_c_U' read by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write6_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~write_back54_U0.hyperedge_size_blk_n) begin
                            if (~hyperedge_size_c855_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c855_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c855_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c855_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c855_U' read by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c855_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back54_U0_U.if_empty_n & write_back54_U0.ap_idle & ~start_for_write_back54_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back54_U0_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0',");
                        end
                    end
                    9: begin
                        if (~write_back54_U0.value_stream_V_V6_blk_n) begin
                            if (~value_stream_6_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_6_V_V_U' written by process 'kernel_pr_kernel_pr.load_value38_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_6_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_6_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_6_V_V_U' read by process 'kernel_pr_kernel_pr.load_value38_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_6_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    19: begin
                        if (ap_done_reg_6 & write_back54_U0.ap_done & ~write_back48_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back48_U0'");
                        end
                    end
                    20: begin
                        if (ap_done_reg_6 & write_back54_U0.ap_done & ~write_back49_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back49_U0'");
                        end
                    end
                    21: begin
                        if (ap_done_reg_6 & write_back54_U0.ap_done & ~write_back50_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back50_U0'");
                        end
                    end
                    22: begin
                        if (ap_done_reg_6 & write_back54_U0.ap_done & ~write_back51_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back51_U0'");
                        end
                    end
                    23: begin
                        if (ap_done_reg_6 & write_back54_U0.ap_done & ~write_back52_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back52_U0'");
                        end
                    end
                    24: begin
                        if (ap_done_reg_6 & write_back54_U0.ap_done & ~write_back53_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back53_U0'");
                        end
                    end
                    26: begin
                        if (ap_done_reg_6 & write_back54_U0.ap_done & ~write_back55_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back55_U0'");
                        end
                    end
                    27: begin
                        if (ap_done_reg_6 & write_back54_U0.ap_done & ~write_back56_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back56_U0'");
                        end
                    end
                    28: begin
                        if (ap_done_reg_6 & write_back54_U0.ap_done & ~write_back57_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back57_U0'");
                        end
                    end
                    29: begin
                        if (ap_done_reg_6 & write_back54_U0.ap_done & ~write_back58_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back58_U0'");
                        end
                    end
                    30: begin
                        if (ap_done_reg_6 & write_back54_U0.ap_done & ~write_back59_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back59_U0'");
                        end
                    end
                    31: begin
                        if (ap_done_reg_6 & write_back54_U0.ap_done & ~write_back60_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back60_U0'");
                        end
                    end
                    32: begin
                        if (ap_done_reg_6 & write_back54_U0.ap_done & ~write_back61_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back61_U0'");
                        end
                    end
                    33: begin
                        if (ap_done_reg_6 & write_back54_U0.ap_done & ~write_back62_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back62_U0'");
                        end
                    end
                    34: begin
                        if (ap_done_reg_6 & write_back54_U0.ap_done & ~write_back63_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back63_U0'");
                        end
                    end
                    endcase
                end
                26 : begin
                    case(index2)
                    0: begin
                        if (~write_back55_U0.H_blk_n) begin
                            if (~H_write7_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write7_c_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write7_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write7_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write7_c_U' read by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write7_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~write_back55_U0.hyperedge_size_blk_n) begin
                            if (~hyperedge_size_c856_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c856_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c856_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c856_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c856_U' read by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c856_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back55_U0_U.if_empty_n & write_back55_U0.ap_idle & ~start_for_write_back55_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back55_U0_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0',");
                        end
                    end
                    10: begin
                        if (~write_back55_U0.value_stream_V_V7_blk_n) begin
                            if (~value_stream_7_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_7_V_V_U' written by process 'kernel_pr_kernel_pr.load_value39_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_7_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_7_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_7_V_V_U' read by process 'kernel_pr_kernel_pr.load_value39_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_7_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    19: begin
                        if (ap_done_reg_7 & write_back55_U0.ap_done & ~write_back48_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back48_U0'");
                        end
                    end
                    20: begin
                        if (ap_done_reg_7 & write_back55_U0.ap_done & ~write_back49_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back49_U0'");
                        end
                    end
                    21: begin
                        if (ap_done_reg_7 & write_back55_U0.ap_done & ~write_back50_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back50_U0'");
                        end
                    end
                    22: begin
                        if (ap_done_reg_7 & write_back55_U0.ap_done & ~write_back51_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back51_U0'");
                        end
                    end
                    23: begin
                        if (ap_done_reg_7 & write_back55_U0.ap_done & ~write_back52_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back52_U0'");
                        end
                    end
                    24: begin
                        if (ap_done_reg_7 & write_back55_U0.ap_done & ~write_back53_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back53_U0'");
                        end
                    end
                    25: begin
                        if (ap_done_reg_7 & write_back55_U0.ap_done & ~write_back54_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back54_U0'");
                        end
                    end
                    27: begin
                        if (ap_done_reg_7 & write_back55_U0.ap_done & ~write_back56_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back56_U0'");
                        end
                    end
                    28: begin
                        if (ap_done_reg_7 & write_back55_U0.ap_done & ~write_back57_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back57_U0'");
                        end
                    end
                    29: begin
                        if (ap_done_reg_7 & write_back55_U0.ap_done & ~write_back58_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back58_U0'");
                        end
                    end
                    30: begin
                        if (ap_done_reg_7 & write_back55_U0.ap_done & ~write_back59_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back59_U0'");
                        end
                    end
                    31: begin
                        if (ap_done_reg_7 & write_back55_U0.ap_done & ~write_back60_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back60_U0'");
                        end
                    end
                    32: begin
                        if (ap_done_reg_7 & write_back55_U0.ap_done & ~write_back61_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back61_U0'");
                        end
                    end
                    33: begin
                        if (ap_done_reg_7 & write_back55_U0.ap_done & ~write_back62_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back62_U0'");
                        end
                    end
                    34: begin
                        if (ap_done_reg_7 & write_back55_U0.ap_done & ~write_back63_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back63_U0'");
                        end
                    end
                    endcase
                end
                27 : begin
                    case(index2)
                    0: begin
                        if (~write_back56_U0.H_blk_n) begin
                            if (~H_write8_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write8_c_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write8_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write8_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write8_c_U' read by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write8_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~write_back56_U0.hyperedge_size_blk_n) begin
                            if (~hyperedge_size_c857_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c857_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c857_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c857_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c857_U' read by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c857_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back56_U0_U.if_empty_n & write_back56_U0.ap_idle & ~start_for_write_back56_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back56_U0_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0',");
                        end
                    end
                    11: begin
                        if (~write_back56_U0.value_stream_V_V8_blk_n) begin
                            if (~value_stream_8_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_8_V_V_U' written by process 'kernel_pr_kernel_pr.load_value40_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_8_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_8_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_8_V_V_U' read by process 'kernel_pr_kernel_pr.load_value40_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_8_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    19: begin
                        if (ap_done_reg_8 & write_back56_U0.ap_done & ~write_back48_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back48_U0'");
                        end
                    end
                    20: begin
                        if (ap_done_reg_8 & write_back56_U0.ap_done & ~write_back49_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back49_U0'");
                        end
                    end
                    21: begin
                        if (ap_done_reg_8 & write_back56_U0.ap_done & ~write_back50_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back50_U0'");
                        end
                    end
                    22: begin
                        if (ap_done_reg_8 & write_back56_U0.ap_done & ~write_back51_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back51_U0'");
                        end
                    end
                    23: begin
                        if (ap_done_reg_8 & write_back56_U0.ap_done & ~write_back52_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back52_U0'");
                        end
                    end
                    24: begin
                        if (ap_done_reg_8 & write_back56_U0.ap_done & ~write_back53_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back53_U0'");
                        end
                    end
                    25: begin
                        if (ap_done_reg_8 & write_back56_U0.ap_done & ~write_back54_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back54_U0'");
                        end
                    end
                    26: begin
                        if (ap_done_reg_8 & write_back56_U0.ap_done & ~write_back55_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back55_U0'");
                        end
                    end
                    28: begin
                        if (ap_done_reg_8 & write_back56_U0.ap_done & ~write_back57_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back57_U0'");
                        end
                    end
                    29: begin
                        if (ap_done_reg_8 & write_back56_U0.ap_done & ~write_back58_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back58_U0'");
                        end
                    end
                    30: begin
                        if (ap_done_reg_8 & write_back56_U0.ap_done & ~write_back59_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back59_U0'");
                        end
                    end
                    31: begin
                        if (ap_done_reg_8 & write_back56_U0.ap_done & ~write_back60_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back60_U0'");
                        end
                    end
                    32: begin
                        if (ap_done_reg_8 & write_back56_U0.ap_done & ~write_back61_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back61_U0'");
                        end
                    end
                    33: begin
                        if (ap_done_reg_8 & write_back56_U0.ap_done & ~write_back62_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back62_U0'");
                        end
                    end
                    34: begin
                        if (ap_done_reg_8 & write_back56_U0.ap_done & ~write_back63_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back63_U0'");
                        end
                    end
                    endcase
                end
                28 : begin
                    case(index2)
                    0: begin
                        if (~write_back57_U0.H_blk_n) begin
                            if (~H_write9_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write9_c_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write9_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write9_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write9_c_U' read by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write9_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~write_back57_U0.hyperedge_size_blk_n) begin
                            if (~hyperedge_size_c858_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c858_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c858_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c858_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c858_U' read by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c858_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back57_U0_U.if_empty_n & write_back57_U0.ap_idle & ~start_for_write_back57_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back57_U0_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0',");
                        end
                    end
                    12: begin
                        if (~write_back57_U0.value_stream_V_V9_blk_n) begin
                            if (~value_stream_9_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_9_V_V_U' written by process 'kernel_pr_kernel_pr.load_value41_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_9_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_9_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_9_V_V_U' read by process 'kernel_pr_kernel_pr.load_value41_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_9_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    19: begin
                        if (ap_done_reg_9 & write_back57_U0.ap_done & ~write_back48_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back48_U0'");
                        end
                    end
                    20: begin
                        if (ap_done_reg_9 & write_back57_U0.ap_done & ~write_back49_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back49_U0'");
                        end
                    end
                    21: begin
                        if (ap_done_reg_9 & write_back57_U0.ap_done & ~write_back50_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back50_U0'");
                        end
                    end
                    22: begin
                        if (ap_done_reg_9 & write_back57_U0.ap_done & ~write_back51_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back51_U0'");
                        end
                    end
                    23: begin
                        if (ap_done_reg_9 & write_back57_U0.ap_done & ~write_back52_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back52_U0'");
                        end
                    end
                    24: begin
                        if (ap_done_reg_9 & write_back57_U0.ap_done & ~write_back53_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back53_U0'");
                        end
                    end
                    25: begin
                        if (ap_done_reg_9 & write_back57_U0.ap_done & ~write_back54_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back54_U0'");
                        end
                    end
                    26: begin
                        if (ap_done_reg_9 & write_back57_U0.ap_done & ~write_back55_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back55_U0'");
                        end
                    end
                    27: begin
                        if (ap_done_reg_9 & write_back57_U0.ap_done & ~write_back56_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back56_U0'");
                        end
                    end
                    29: begin
                        if (ap_done_reg_9 & write_back57_U0.ap_done & ~write_back58_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back58_U0'");
                        end
                    end
                    30: begin
                        if (ap_done_reg_9 & write_back57_U0.ap_done & ~write_back59_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back59_U0'");
                        end
                    end
                    31: begin
                        if (ap_done_reg_9 & write_back57_U0.ap_done & ~write_back60_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back60_U0'");
                        end
                    end
                    32: begin
                        if (ap_done_reg_9 & write_back57_U0.ap_done & ~write_back61_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back61_U0'");
                        end
                    end
                    33: begin
                        if (ap_done_reg_9 & write_back57_U0.ap_done & ~write_back62_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back62_U0'");
                        end
                    end
                    34: begin
                        if (ap_done_reg_9 & write_back57_U0.ap_done & ~write_back63_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back63_U0'");
                        end
                    end
                    endcase
                end
                29 : begin
                    case(index2)
                    0: begin
                        if (~write_back58_U0.H_blk_n) begin
                            if (~H_write10_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write10_c_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write10_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write10_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write10_c_U' read by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write10_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~write_back58_U0.hyperedge_size_blk_n) begin
                            if (~hyperedge_size_c859_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c859_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c859_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c859_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c859_U' read by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c859_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back58_U0_U.if_empty_n & write_back58_U0.ap_idle & ~start_for_write_back58_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back58_U0_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0',");
                        end
                    end
                    13: begin
                        if (~write_back58_U0.value_stream_V_V10_blk_n) begin
                            if (~value_stream_10_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_10_V_V_U' written by process 'kernel_pr_kernel_pr.load_value42_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_10_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_10_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_10_V_V_U' read by process 'kernel_pr_kernel_pr.load_value42_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_10_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    19: begin
                        if (ap_done_reg_10 & write_back58_U0.ap_done & ~write_back48_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back48_U0'");
                        end
                    end
                    20: begin
                        if (ap_done_reg_10 & write_back58_U0.ap_done & ~write_back49_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back49_U0'");
                        end
                    end
                    21: begin
                        if (ap_done_reg_10 & write_back58_U0.ap_done & ~write_back50_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back50_U0'");
                        end
                    end
                    22: begin
                        if (ap_done_reg_10 & write_back58_U0.ap_done & ~write_back51_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back51_U0'");
                        end
                    end
                    23: begin
                        if (ap_done_reg_10 & write_back58_U0.ap_done & ~write_back52_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back52_U0'");
                        end
                    end
                    24: begin
                        if (ap_done_reg_10 & write_back58_U0.ap_done & ~write_back53_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back53_U0'");
                        end
                    end
                    25: begin
                        if (ap_done_reg_10 & write_back58_U0.ap_done & ~write_back54_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back54_U0'");
                        end
                    end
                    26: begin
                        if (ap_done_reg_10 & write_back58_U0.ap_done & ~write_back55_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back55_U0'");
                        end
                    end
                    27: begin
                        if (ap_done_reg_10 & write_back58_U0.ap_done & ~write_back56_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back56_U0'");
                        end
                    end
                    28: begin
                        if (ap_done_reg_10 & write_back58_U0.ap_done & ~write_back57_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back57_U0'");
                        end
                    end
                    30: begin
                        if (ap_done_reg_10 & write_back58_U0.ap_done & ~write_back59_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back59_U0'");
                        end
                    end
                    31: begin
                        if (ap_done_reg_10 & write_back58_U0.ap_done & ~write_back60_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back60_U0'");
                        end
                    end
                    32: begin
                        if (ap_done_reg_10 & write_back58_U0.ap_done & ~write_back61_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back61_U0'");
                        end
                    end
                    33: begin
                        if (ap_done_reg_10 & write_back58_U0.ap_done & ~write_back62_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back62_U0'");
                        end
                    end
                    34: begin
                        if (ap_done_reg_10 & write_back58_U0.ap_done & ~write_back63_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back63_U0'");
                        end
                    end
                    endcase
                end
                30 : begin
                    case(index2)
                    0: begin
                        if (~write_back59_U0.H_blk_n) begin
                            if (~H_write11_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write11_c_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write11_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write11_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write11_c_U' read by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write11_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~write_back59_U0.hyperedge_size_blk_n) begin
                            if (~hyperedge_size_c860_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c860_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c860_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c860_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c860_U' read by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c860_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back59_U0_U.if_empty_n & write_back59_U0.ap_idle & ~start_for_write_back59_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back59_U0_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0',");
                        end
                    end
                    14: begin
                        if (~write_back59_U0.value_stream_V_V11_blk_n) begin
                            if (~value_stream_11_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_11_V_V_U' written by process 'kernel_pr_kernel_pr.load_value43_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_11_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_11_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_11_V_V_U' read by process 'kernel_pr_kernel_pr.load_value43_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_11_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    19: begin
                        if (ap_done_reg_11 & write_back59_U0.ap_done & ~write_back48_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back48_U0'");
                        end
                    end
                    20: begin
                        if (ap_done_reg_11 & write_back59_U0.ap_done & ~write_back49_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back49_U0'");
                        end
                    end
                    21: begin
                        if (ap_done_reg_11 & write_back59_U0.ap_done & ~write_back50_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back50_U0'");
                        end
                    end
                    22: begin
                        if (ap_done_reg_11 & write_back59_U0.ap_done & ~write_back51_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back51_U0'");
                        end
                    end
                    23: begin
                        if (ap_done_reg_11 & write_back59_U0.ap_done & ~write_back52_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back52_U0'");
                        end
                    end
                    24: begin
                        if (ap_done_reg_11 & write_back59_U0.ap_done & ~write_back53_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back53_U0'");
                        end
                    end
                    25: begin
                        if (ap_done_reg_11 & write_back59_U0.ap_done & ~write_back54_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back54_U0'");
                        end
                    end
                    26: begin
                        if (ap_done_reg_11 & write_back59_U0.ap_done & ~write_back55_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back55_U0'");
                        end
                    end
                    27: begin
                        if (ap_done_reg_11 & write_back59_U0.ap_done & ~write_back56_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back56_U0'");
                        end
                    end
                    28: begin
                        if (ap_done_reg_11 & write_back59_U0.ap_done & ~write_back57_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back57_U0'");
                        end
                    end
                    29: begin
                        if (ap_done_reg_11 & write_back59_U0.ap_done & ~write_back58_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back58_U0'");
                        end
                    end
                    31: begin
                        if (ap_done_reg_11 & write_back59_U0.ap_done & ~write_back60_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back60_U0'");
                        end
                    end
                    32: begin
                        if (ap_done_reg_11 & write_back59_U0.ap_done & ~write_back61_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back61_U0'");
                        end
                    end
                    33: begin
                        if (ap_done_reg_11 & write_back59_U0.ap_done & ~write_back62_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back62_U0'");
                        end
                    end
                    34: begin
                        if (ap_done_reg_11 & write_back59_U0.ap_done & ~write_back63_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back63_U0'");
                        end
                    end
                    endcase
                end
                31 : begin
                    case(index2)
                    0: begin
                        if (~write_back60_U0.H_blk_n) begin
                            if (~H_write12_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write12_c_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write12_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write12_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write12_c_U' read by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write12_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~write_back60_U0.hyperedge_size_blk_n) begin
                            if (~hyperedge_size_c861_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c861_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c861_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c861_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c861_U' read by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c861_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back60_U0_U.if_empty_n & write_back60_U0.ap_idle & ~start_for_write_back60_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back60_U0_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0',");
                        end
                    end
                    15: begin
                        if (~write_back60_U0.value_stream_V_V12_blk_n) begin
                            if (~value_stream_12_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_12_V_V_U' written by process 'kernel_pr_kernel_pr.load_value44_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_12_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_12_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_12_V_V_U' read by process 'kernel_pr_kernel_pr.load_value44_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_12_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    19: begin
                        if (ap_done_reg_12 & write_back60_U0.ap_done & ~write_back48_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back48_U0'");
                        end
                    end
                    20: begin
                        if (ap_done_reg_12 & write_back60_U0.ap_done & ~write_back49_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back49_U0'");
                        end
                    end
                    21: begin
                        if (ap_done_reg_12 & write_back60_U0.ap_done & ~write_back50_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back50_U0'");
                        end
                    end
                    22: begin
                        if (ap_done_reg_12 & write_back60_U0.ap_done & ~write_back51_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back51_U0'");
                        end
                    end
                    23: begin
                        if (ap_done_reg_12 & write_back60_U0.ap_done & ~write_back52_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back52_U0'");
                        end
                    end
                    24: begin
                        if (ap_done_reg_12 & write_back60_U0.ap_done & ~write_back53_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back53_U0'");
                        end
                    end
                    25: begin
                        if (ap_done_reg_12 & write_back60_U0.ap_done & ~write_back54_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back54_U0'");
                        end
                    end
                    26: begin
                        if (ap_done_reg_12 & write_back60_U0.ap_done & ~write_back55_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back55_U0'");
                        end
                    end
                    27: begin
                        if (ap_done_reg_12 & write_back60_U0.ap_done & ~write_back56_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back56_U0'");
                        end
                    end
                    28: begin
                        if (ap_done_reg_12 & write_back60_U0.ap_done & ~write_back57_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back57_U0'");
                        end
                    end
                    29: begin
                        if (ap_done_reg_12 & write_back60_U0.ap_done & ~write_back58_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back58_U0'");
                        end
                    end
                    30: begin
                        if (ap_done_reg_12 & write_back60_U0.ap_done & ~write_back59_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back59_U0'");
                        end
                    end
                    32: begin
                        if (ap_done_reg_12 & write_back60_U0.ap_done & ~write_back61_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back61_U0'");
                        end
                    end
                    33: begin
                        if (ap_done_reg_12 & write_back60_U0.ap_done & ~write_back62_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back62_U0'");
                        end
                    end
                    34: begin
                        if (ap_done_reg_12 & write_back60_U0.ap_done & ~write_back63_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back63_U0'");
                        end
                    end
                    endcase
                end
                32 : begin
                    case(index2)
                    0: begin
                        if (~write_back61_U0.H_blk_n) begin
                            if (~H_write13_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write13_c_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write13_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write13_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write13_c_U' read by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write13_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~write_back61_U0.hyperedge_size_blk_n) begin
                            if (~hyperedge_size_c862_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c862_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c862_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c862_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c862_U' read by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c862_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back61_U0_U.if_empty_n & write_back61_U0.ap_idle & ~start_for_write_back61_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back61_U0_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0',");
                        end
                    end
                    16: begin
                        if (~write_back61_U0.value_stream_V_V13_blk_n) begin
                            if (~value_stream_13_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_13_V_V_U' written by process 'kernel_pr_kernel_pr.load_value45_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_13_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_13_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_13_V_V_U' read by process 'kernel_pr_kernel_pr.load_value45_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_13_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    19: begin
                        if (ap_done_reg_13 & write_back61_U0.ap_done & ~write_back48_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back48_U0'");
                        end
                    end
                    20: begin
                        if (ap_done_reg_13 & write_back61_U0.ap_done & ~write_back49_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back49_U0'");
                        end
                    end
                    21: begin
                        if (ap_done_reg_13 & write_back61_U0.ap_done & ~write_back50_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back50_U0'");
                        end
                    end
                    22: begin
                        if (ap_done_reg_13 & write_back61_U0.ap_done & ~write_back51_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back51_U0'");
                        end
                    end
                    23: begin
                        if (ap_done_reg_13 & write_back61_U0.ap_done & ~write_back52_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back52_U0'");
                        end
                    end
                    24: begin
                        if (ap_done_reg_13 & write_back61_U0.ap_done & ~write_back53_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back53_U0'");
                        end
                    end
                    25: begin
                        if (ap_done_reg_13 & write_back61_U0.ap_done & ~write_back54_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back54_U0'");
                        end
                    end
                    26: begin
                        if (ap_done_reg_13 & write_back61_U0.ap_done & ~write_back55_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back55_U0'");
                        end
                    end
                    27: begin
                        if (ap_done_reg_13 & write_back61_U0.ap_done & ~write_back56_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back56_U0'");
                        end
                    end
                    28: begin
                        if (ap_done_reg_13 & write_back61_U0.ap_done & ~write_back57_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back57_U0'");
                        end
                    end
                    29: begin
                        if (ap_done_reg_13 & write_back61_U0.ap_done & ~write_back58_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back58_U0'");
                        end
                    end
                    30: begin
                        if (ap_done_reg_13 & write_back61_U0.ap_done & ~write_back59_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back59_U0'");
                        end
                    end
                    31: begin
                        if (ap_done_reg_13 & write_back61_U0.ap_done & ~write_back60_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back60_U0'");
                        end
                    end
                    33: begin
                        if (ap_done_reg_13 & write_back61_U0.ap_done & ~write_back62_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back62_U0'");
                        end
                    end
                    34: begin
                        if (ap_done_reg_13 & write_back61_U0.ap_done & ~write_back63_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back63_U0'");
                        end
                    end
                    endcase
                end
                33 : begin
                    case(index2)
                    0: begin
                        if (~write_back62_U0.H_blk_n) begin
                            if (~H_write14_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write14_c_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write14_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write14_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write14_c_U' read by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write14_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~write_back62_U0.hyperedge_size_blk_n) begin
                            if (~hyperedge_size_c863_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c863_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c863_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c863_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c863_U' read by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c863_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back62_U0_U.if_empty_n & write_back62_U0.ap_idle & ~start_for_write_back62_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back62_U0_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0',");
                        end
                    end
                    17: begin
                        if (~write_back62_U0.value_stream_V_V14_blk_n) begin
                            if (~value_stream_14_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_14_V_V_U' written by process 'kernel_pr_kernel_pr.load_value46_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_14_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_14_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_14_V_V_U' read by process 'kernel_pr_kernel_pr.load_value46_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_14_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    19: begin
                        if (ap_done_reg_14 & write_back62_U0.ap_done & ~write_back48_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back48_U0'");
                        end
                    end
                    20: begin
                        if (ap_done_reg_14 & write_back62_U0.ap_done & ~write_back49_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back49_U0'");
                        end
                    end
                    21: begin
                        if (ap_done_reg_14 & write_back62_U0.ap_done & ~write_back50_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back50_U0'");
                        end
                    end
                    22: begin
                        if (ap_done_reg_14 & write_back62_U0.ap_done & ~write_back51_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back51_U0'");
                        end
                    end
                    23: begin
                        if (ap_done_reg_14 & write_back62_U0.ap_done & ~write_back52_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back52_U0'");
                        end
                    end
                    24: begin
                        if (ap_done_reg_14 & write_back62_U0.ap_done & ~write_back53_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back53_U0'");
                        end
                    end
                    25: begin
                        if (ap_done_reg_14 & write_back62_U0.ap_done & ~write_back54_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back54_U0'");
                        end
                    end
                    26: begin
                        if (ap_done_reg_14 & write_back62_U0.ap_done & ~write_back55_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back55_U0'");
                        end
                    end
                    27: begin
                        if (ap_done_reg_14 & write_back62_U0.ap_done & ~write_back56_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back56_U0'");
                        end
                    end
                    28: begin
                        if (ap_done_reg_14 & write_back62_U0.ap_done & ~write_back57_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back57_U0'");
                        end
                    end
                    29: begin
                        if (ap_done_reg_14 & write_back62_U0.ap_done & ~write_back58_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back58_U0'");
                        end
                    end
                    30: begin
                        if (ap_done_reg_14 & write_back62_U0.ap_done & ~write_back59_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back59_U0'");
                        end
                    end
                    31: begin
                        if (ap_done_reg_14 & write_back62_U0.ap_done & ~write_back60_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back60_U0'");
                        end
                    end
                    32: begin
                        if (ap_done_reg_14 & write_back62_U0.ap_done & ~write_back61_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back61_U0'");
                        end
                    end
                    34: begin
                        if (ap_done_reg_14 & write_back62_U0.ap_done & ~write_back63_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back63_U0'");
                        end
                    end
                    endcase
                end
                34 : begin
                    case(index2)
                    0: begin
                        if (~write_back63_U0.H_blk_n) begin
                            if (~H_write15_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.H_write15_c_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write15_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~H_write15_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.H_write15_c_U' read by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.H_write15_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~write_back63_U0.hyperedge_size_blk_n) begin
                            if (~hyperedge_size_c864_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.hyperedge_size_c864_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c864_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~hyperedge_size_c864_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.hyperedge_size_c864_U' read by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.hyperedge_size_c864_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~start_for_write_back63_U0_U.if_empty_n & write_back63_U0.ap_idle & ~start_for_write_back63_U0_U.if_write) begin
                            $display("//      Blocked by missing 'ap_start' from start propagation FIFO 'kernel_pr_kernel_pr.start_for_write_back63_U0_U' written by process 'kernel_pr_kernel_pr.kernel_pr_entry98_U0',");
                        end
                    end
                    18: begin
                        if (~write_back63_U0.value_stream_V_V15_blk_n) begin
                            if (~value_stream_15_V_V_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'kernel_pr_kernel_pr.value_stream_15_V_V_U' written by process 'kernel_pr_kernel_pr.load_value47_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_15_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~value_stream_15_V_V_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'kernel_pr_kernel_pr.value_stream_15_V_V_U' read by process 'kernel_pr_kernel_pr.load_value47_U0'");
                                $fdisplay(fp, "Dependence_Channel_path kernel_pr_kernel_pr.value_stream_15_V_V_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    19: begin
                        if (ap_done_reg_15 & write_back63_U0.ap_done & ~write_back48_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back48_U0'");
                        end
                    end
                    20: begin
                        if (ap_done_reg_15 & write_back63_U0.ap_done & ~write_back49_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back49_U0'");
                        end
                    end
                    21: begin
                        if (ap_done_reg_15 & write_back63_U0.ap_done & ~write_back50_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back50_U0'");
                        end
                    end
                    22: begin
                        if (ap_done_reg_15 & write_back63_U0.ap_done & ~write_back51_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back51_U0'");
                        end
                    end
                    23: begin
                        if (ap_done_reg_15 & write_back63_U0.ap_done & ~write_back52_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back52_U0'");
                        end
                    end
                    24: begin
                        if (ap_done_reg_15 & write_back63_U0.ap_done & ~write_back53_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back53_U0'");
                        end
                    end
                    25: begin
                        if (ap_done_reg_15 & write_back63_U0.ap_done & ~write_back54_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back54_U0'");
                        end
                    end
                    26: begin
                        if (ap_done_reg_15 & write_back63_U0.ap_done & ~write_back55_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back55_U0'");
                        end
                    end
                    27: begin
                        if (ap_done_reg_15 & write_back63_U0.ap_done & ~write_back56_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back56_U0'");
                        end
                    end
                    28: begin
                        if (ap_done_reg_15 & write_back63_U0.ap_done & ~write_back57_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back57_U0'");
                        end
                    end
                    29: begin
                        if (ap_done_reg_15 & write_back63_U0.ap_done & ~write_back58_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back58_U0'");
                        end
                    end
                    30: begin
                        if (ap_done_reg_15 & write_back63_U0.ap_done & ~write_back59_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back59_U0'");
                        end
                    end
                    31: begin
                        if (ap_done_reg_15 & write_back63_U0.ap_done & ~write_back60_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back60_U0'");
                        end
                    end
                    32: begin
                        if (ap_done_reg_15 & write_back63_U0.ap_done & ~write_back61_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back61_U0'");
                        end
                    end
                    33: begin
                        if (ap_done_reg_15 & write_back63_U0.ap_done & ~write_back62_U0.ap_done) begin
                            $display("//      Blocked by output sync logic with process : 'kernel_pr_kernel_pr.write_back62_U0'");
                        end
                    end
                    endcase
                end
            endcase
        end
    endtask

    // report
    initial begin : report_deadlock
        integer cycle_id;
        integer cycle_comp_id;
        integer record_time;
        wait (reset == 1);
        cycle_id = 1;
        record_time = 0;
        while (1) begin
            @ (negedge clock);
            case (CS_fsm)
                ST_DL_DETECTED: begin
                    cycle_comp_id = 2;
                    if (dl_detect_reg != dl_done_reg) begin
                        if (dl_done_reg == 'b0) begin
                            print_dl_head;
                            record_time = $time;
                        end
                        print_cycle_start(proc_path(origin), cycle_id);
                        cycle_id = cycle_id + 1;
                    end
                    else begin
                        print_dl_end((cycle_id - 1),record_time);
                        find_df_deadlock = 1;
                        @(negedge clock);
                        $finish;
                    end
                end
                ST_DL_REPORT: begin
                    if ((|(dl_in_vec)) & ~(|(dl_in_vec & origin_reg))) begin
                        print_cycle_chan_comp(dl_in_vec_reg, dl_in_vec);
                        print_cycle_proc_comp(proc_path(dl_in_vec), cycle_comp_id);
                        cycle_comp_id = cycle_comp_id + 1;
                    end
                    else begin
                        print_cycle_chan_comp(dl_in_vec_reg, dl_in_vec);
                    end
                end
            endcase
        end
    end
 
