
    wire reset;
    wire clock;
    assign reset = ap_rst_n;
    assign clock = ap_clk;
    wire [33:0] proc_0_data_FIFO_blk;
    wire [33:0] proc_0_data_PIPO_blk;
    wire [33:0] proc_0_start_FIFO_blk;
    wire [33:0] proc_0_TLF_FIFO_blk;
    wire [33:0] proc_0_input_sync_blk;
    wire [33:0] proc_0_output_sync_blk;
    wire [33:0] proc_dep_vld_vec_0;
    reg [33:0] proc_dep_vld_vec_0_reg;
    wire [33:0] in_chan_dep_vld_vec_0;
    wire [1189:0] in_chan_dep_data_vec_0;
    wire [33:0] token_in_vec_0;
    wire [33:0] out_chan_dep_vld_vec_0;
    wire [34:0] out_chan_dep_data_0;
    wire [33:0] token_out_vec_0;
    wire dl_detect_out_0;
    wire dep_chan_vld_1_0;
    wire [34:0] dep_chan_data_1_0;
    wire token_1_0;
    wire dep_chan_vld_2_0;
    wire [34:0] dep_chan_data_2_0;
    wire token_2_0;
    wire dep_chan_vld_3_0;
    wire [34:0] dep_chan_data_3_0;
    wire token_3_0;
    wire dep_chan_vld_4_0;
    wire [34:0] dep_chan_data_4_0;
    wire token_4_0;
    wire dep_chan_vld_5_0;
    wire [34:0] dep_chan_data_5_0;
    wire token_5_0;
    wire dep_chan_vld_6_0;
    wire [34:0] dep_chan_data_6_0;
    wire token_6_0;
    wire dep_chan_vld_7_0;
    wire [34:0] dep_chan_data_7_0;
    wire token_7_0;
    wire dep_chan_vld_8_0;
    wire [34:0] dep_chan_data_8_0;
    wire token_8_0;
    wire dep_chan_vld_9_0;
    wire [34:0] dep_chan_data_9_0;
    wire token_9_0;
    wire dep_chan_vld_10_0;
    wire [34:0] dep_chan_data_10_0;
    wire token_10_0;
    wire dep_chan_vld_11_0;
    wire [34:0] dep_chan_data_11_0;
    wire token_11_0;
    wire dep_chan_vld_12_0;
    wire [34:0] dep_chan_data_12_0;
    wire token_12_0;
    wire dep_chan_vld_13_0;
    wire [34:0] dep_chan_data_13_0;
    wire token_13_0;
    wire dep_chan_vld_14_0;
    wire [34:0] dep_chan_data_14_0;
    wire token_14_0;
    wire dep_chan_vld_15_0;
    wire [34:0] dep_chan_data_15_0;
    wire token_15_0;
    wire dep_chan_vld_16_0;
    wire [34:0] dep_chan_data_16_0;
    wire token_16_0;
    wire dep_chan_vld_17_0;
    wire [34:0] dep_chan_data_17_0;
    wire token_17_0;
    wire dep_chan_vld_18_0;
    wire [34:0] dep_chan_data_18_0;
    wire token_18_0;
    wire dep_chan_vld_19_0;
    wire [34:0] dep_chan_data_19_0;
    wire token_19_0;
    wire dep_chan_vld_20_0;
    wire [34:0] dep_chan_data_20_0;
    wire token_20_0;
    wire dep_chan_vld_21_0;
    wire [34:0] dep_chan_data_21_0;
    wire token_21_0;
    wire dep_chan_vld_22_0;
    wire [34:0] dep_chan_data_22_0;
    wire token_22_0;
    wire dep_chan_vld_23_0;
    wire [34:0] dep_chan_data_23_0;
    wire token_23_0;
    wire dep_chan_vld_24_0;
    wire [34:0] dep_chan_data_24_0;
    wire token_24_0;
    wire dep_chan_vld_25_0;
    wire [34:0] dep_chan_data_25_0;
    wire token_25_0;
    wire dep_chan_vld_26_0;
    wire [34:0] dep_chan_data_26_0;
    wire token_26_0;
    wire dep_chan_vld_27_0;
    wire [34:0] dep_chan_data_27_0;
    wire token_27_0;
    wire dep_chan_vld_28_0;
    wire [34:0] dep_chan_data_28_0;
    wire token_28_0;
    wire dep_chan_vld_29_0;
    wire [34:0] dep_chan_data_29_0;
    wire token_29_0;
    wire dep_chan_vld_30_0;
    wire [34:0] dep_chan_data_30_0;
    wire token_30_0;
    wire dep_chan_vld_31_0;
    wire [34:0] dep_chan_data_31_0;
    wire token_31_0;
    wire dep_chan_vld_32_0;
    wire [34:0] dep_chan_data_32_0;
    wire token_32_0;
    wire dep_chan_vld_33_0;
    wire [34:0] dep_chan_data_33_0;
    wire token_33_0;
    wire dep_chan_vld_34_0;
    wire [34:0] dep_chan_data_34_0;
    wire token_34_0;
    wire [17:0] proc_1_data_FIFO_blk;
    wire [17:0] proc_1_data_PIPO_blk;
    wire [17:0] proc_1_start_FIFO_blk;
    wire [17:0] proc_1_TLF_FIFO_blk;
    wire [17:0] proc_1_input_sync_blk;
    wire [17:0] proc_1_output_sync_blk;
    wire [17:0] proc_dep_vld_vec_1;
    reg [17:0] proc_dep_vld_vec_1_reg;
    wire [17:0] in_chan_dep_vld_vec_1;
    wire [629:0] in_chan_dep_data_vec_1;
    wire [17:0] token_in_vec_1;
    wire [17:0] out_chan_dep_vld_vec_1;
    wire [34:0] out_chan_dep_data_1;
    wire [17:0] token_out_vec_1;
    wire dl_detect_out_1;
    wire dep_chan_vld_0_1;
    wire [34:0] dep_chan_data_0_1;
    wire token_0_1;
    wire dep_chan_vld_2_1;
    wire [34:0] dep_chan_data_2_1;
    wire token_2_1;
    wire dep_chan_vld_3_1;
    wire [34:0] dep_chan_data_3_1;
    wire token_3_1;
    wire dep_chan_vld_4_1;
    wire [34:0] dep_chan_data_4_1;
    wire token_4_1;
    wire dep_chan_vld_5_1;
    wire [34:0] dep_chan_data_5_1;
    wire token_5_1;
    wire dep_chan_vld_6_1;
    wire [34:0] dep_chan_data_6_1;
    wire token_6_1;
    wire dep_chan_vld_7_1;
    wire [34:0] dep_chan_data_7_1;
    wire token_7_1;
    wire dep_chan_vld_8_1;
    wire [34:0] dep_chan_data_8_1;
    wire token_8_1;
    wire dep_chan_vld_9_1;
    wire [34:0] dep_chan_data_9_1;
    wire token_9_1;
    wire dep_chan_vld_10_1;
    wire [34:0] dep_chan_data_10_1;
    wire token_10_1;
    wire dep_chan_vld_11_1;
    wire [34:0] dep_chan_data_11_1;
    wire token_11_1;
    wire dep_chan_vld_12_1;
    wire [34:0] dep_chan_data_12_1;
    wire token_12_1;
    wire dep_chan_vld_13_1;
    wire [34:0] dep_chan_data_13_1;
    wire token_13_1;
    wire dep_chan_vld_14_1;
    wire [34:0] dep_chan_data_14_1;
    wire token_14_1;
    wire dep_chan_vld_15_1;
    wire [34:0] dep_chan_data_15_1;
    wire token_15_1;
    wire dep_chan_vld_16_1;
    wire [34:0] dep_chan_data_16_1;
    wire token_16_1;
    wire dep_chan_vld_17_1;
    wire [34:0] dep_chan_data_17_1;
    wire token_17_1;
    wire dep_chan_vld_18_1;
    wire [34:0] dep_chan_data_18_1;
    wire token_18_1;
    wire [17:0] proc_2_data_FIFO_blk;
    wire [17:0] proc_2_data_PIPO_blk;
    wire [17:0] proc_2_start_FIFO_blk;
    wire [17:0] proc_2_TLF_FIFO_blk;
    wire [17:0] proc_2_input_sync_blk;
    wire [17:0] proc_2_output_sync_blk;
    wire [17:0] proc_dep_vld_vec_2;
    reg [17:0] proc_dep_vld_vec_2_reg;
    wire [17:0] in_chan_dep_vld_vec_2;
    wire [629:0] in_chan_dep_data_vec_2;
    wire [17:0] token_in_vec_2;
    wire [17:0] out_chan_dep_vld_vec_2;
    wire [34:0] out_chan_dep_data_2;
    wire [17:0] token_out_vec_2;
    wire dl_detect_out_2;
    wire dep_chan_vld_0_2;
    wire [34:0] dep_chan_data_0_2;
    wire token_0_2;
    wire dep_chan_vld_1_2;
    wire [34:0] dep_chan_data_1_2;
    wire token_1_2;
    wire dep_chan_vld_3_2;
    wire [34:0] dep_chan_data_3_2;
    wire token_3_2;
    wire dep_chan_vld_4_2;
    wire [34:0] dep_chan_data_4_2;
    wire token_4_2;
    wire dep_chan_vld_5_2;
    wire [34:0] dep_chan_data_5_2;
    wire token_5_2;
    wire dep_chan_vld_6_2;
    wire [34:0] dep_chan_data_6_2;
    wire token_6_2;
    wire dep_chan_vld_7_2;
    wire [34:0] dep_chan_data_7_2;
    wire token_7_2;
    wire dep_chan_vld_8_2;
    wire [34:0] dep_chan_data_8_2;
    wire token_8_2;
    wire dep_chan_vld_9_2;
    wire [34:0] dep_chan_data_9_2;
    wire token_9_2;
    wire dep_chan_vld_10_2;
    wire [34:0] dep_chan_data_10_2;
    wire token_10_2;
    wire dep_chan_vld_11_2;
    wire [34:0] dep_chan_data_11_2;
    wire token_11_2;
    wire dep_chan_vld_12_2;
    wire [34:0] dep_chan_data_12_2;
    wire token_12_2;
    wire dep_chan_vld_13_2;
    wire [34:0] dep_chan_data_13_2;
    wire token_13_2;
    wire dep_chan_vld_14_2;
    wire [34:0] dep_chan_data_14_2;
    wire token_14_2;
    wire dep_chan_vld_15_2;
    wire [34:0] dep_chan_data_15_2;
    wire token_15_2;
    wire dep_chan_vld_16_2;
    wire [34:0] dep_chan_data_16_2;
    wire token_16_2;
    wire dep_chan_vld_17_2;
    wire [34:0] dep_chan_data_17_2;
    wire token_17_2;
    wire dep_chan_vld_18_2;
    wire [34:0] dep_chan_data_18_2;
    wire token_18_2;
    wire [18:0] proc_3_data_FIFO_blk;
    wire [18:0] proc_3_data_PIPO_blk;
    wire [18:0] proc_3_start_FIFO_blk;
    wire [18:0] proc_3_TLF_FIFO_blk;
    wire [18:0] proc_3_input_sync_blk;
    wire [18:0] proc_3_output_sync_blk;
    wire [18:0] proc_dep_vld_vec_3;
    reg [18:0] proc_dep_vld_vec_3_reg;
    wire [18:0] in_chan_dep_vld_vec_3;
    wire [664:0] in_chan_dep_data_vec_3;
    wire [18:0] token_in_vec_3;
    wire [18:0] out_chan_dep_vld_vec_3;
    wire [34:0] out_chan_dep_data_3;
    wire [18:0] token_out_vec_3;
    wire dl_detect_out_3;
    wire dep_chan_vld_0_3;
    wire [34:0] dep_chan_data_0_3;
    wire token_0_3;
    wire dep_chan_vld_1_3;
    wire [34:0] dep_chan_data_1_3;
    wire token_1_3;
    wire dep_chan_vld_2_3;
    wire [34:0] dep_chan_data_2_3;
    wire token_2_3;
    wire dep_chan_vld_4_3;
    wire [34:0] dep_chan_data_4_3;
    wire token_4_3;
    wire dep_chan_vld_5_3;
    wire [34:0] dep_chan_data_5_3;
    wire token_5_3;
    wire dep_chan_vld_6_3;
    wire [34:0] dep_chan_data_6_3;
    wire token_6_3;
    wire dep_chan_vld_7_3;
    wire [34:0] dep_chan_data_7_3;
    wire token_7_3;
    wire dep_chan_vld_8_3;
    wire [34:0] dep_chan_data_8_3;
    wire token_8_3;
    wire dep_chan_vld_9_3;
    wire [34:0] dep_chan_data_9_3;
    wire token_9_3;
    wire dep_chan_vld_10_3;
    wire [34:0] dep_chan_data_10_3;
    wire token_10_3;
    wire dep_chan_vld_11_3;
    wire [34:0] dep_chan_data_11_3;
    wire token_11_3;
    wire dep_chan_vld_12_3;
    wire [34:0] dep_chan_data_12_3;
    wire token_12_3;
    wire dep_chan_vld_13_3;
    wire [34:0] dep_chan_data_13_3;
    wire token_13_3;
    wire dep_chan_vld_14_3;
    wire [34:0] dep_chan_data_14_3;
    wire token_14_3;
    wire dep_chan_vld_15_3;
    wire [34:0] dep_chan_data_15_3;
    wire token_15_3;
    wire dep_chan_vld_16_3;
    wire [34:0] dep_chan_data_16_3;
    wire token_16_3;
    wire dep_chan_vld_17_3;
    wire [34:0] dep_chan_data_17_3;
    wire token_17_3;
    wire dep_chan_vld_18_3;
    wire [34:0] dep_chan_data_18_3;
    wire token_18_3;
    wire dep_chan_vld_19_3;
    wire [34:0] dep_chan_data_19_3;
    wire token_19_3;
    wire [18:0] proc_4_data_FIFO_blk;
    wire [18:0] proc_4_data_PIPO_blk;
    wire [18:0] proc_4_start_FIFO_blk;
    wire [18:0] proc_4_TLF_FIFO_blk;
    wire [18:0] proc_4_input_sync_blk;
    wire [18:0] proc_4_output_sync_blk;
    wire [18:0] proc_dep_vld_vec_4;
    reg [18:0] proc_dep_vld_vec_4_reg;
    wire [18:0] in_chan_dep_vld_vec_4;
    wire [664:0] in_chan_dep_data_vec_4;
    wire [18:0] token_in_vec_4;
    wire [18:0] out_chan_dep_vld_vec_4;
    wire [34:0] out_chan_dep_data_4;
    wire [18:0] token_out_vec_4;
    wire dl_detect_out_4;
    wire dep_chan_vld_0_4;
    wire [34:0] dep_chan_data_0_4;
    wire token_0_4;
    wire dep_chan_vld_1_4;
    wire [34:0] dep_chan_data_1_4;
    wire token_1_4;
    wire dep_chan_vld_2_4;
    wire [34:0] dep_chan_data_2_4;
    wire token_2_4;
    wire dep_chan_vld_3_4;
    wire [34:0] dep_chan_data_3_4;
    wire token_3_4;
    wire dep_chan_vld_5_4;
    wire [34:0] dep_chan_data_5_4;
    wire token_5_4;
    wire dep_chan_vld_6_4;
    wire [34:0] dep_chan_data_6_4;
    wire token_6_4;
    wire dep_chan_vld_7_4;
    wire [34:0] dep_chan_data_7_4;
    wire token_7_4;
    wire dep_chan_vld_8_4;
    wire [34:0] dep_chan_data_8_4;
    wire token_8_4;
    wire dep_chan_vld_9_4;
    wire [34:0] dep_chan_data_9_4;
    wire token_9_4;
    wire dep_chan_vld_10_4;
    wire [34:0] dep_chan_data_10_4;
    wire token_10_4;
    wire dep_chan_vld_11_4;
    wire [34:0] dep_chan_data_11_4;
    wire token_11_4;
    wire dep_chan_vld_12_4;
    wire [34:0] dep_chan_data_12_4;
    wire token_12_4;
    wire dep_chan_vld_13_4;
    wire [34:0] dep_chan_data_13_4;
    wire token_13_4;
    wire dep_chan_vld_14_4;
    wire [34:0] dep_chan_data_14_4;
    wire token_14_4;
    wire dep_chan_vld_15_4;
    wire [34:0] dep_chan_data_15_4;
    wire token_15_4;
    wire dep_chan_vld_16_4;
    wire [34:0] dep_chan_data_16_4;
    wire token_16_4;
    wire dep_chan_vld_17_4;
    wire [34:0] dep_chan_data_17_4;
    wire token_17_4;
    wire dep_chan_vld_18_4;
    wire [34:0] dep_chan_data_18_4;
    wire token_18_4;
    wire dep_chan_vld_20_4;
    wire [34:0] dep_chan_data_20_4;
    wire token_20_4;
    wire [18:0] proc_5_data_FIFO_blk;
    wire [18:0] proc_5_data_PIPO_blk;
    wire [18:0] proc_5_start_FIFO_blk;
    wire [18:0] proc_5_TLF_FIFO_blk;
    wire [18:0] proc_5_input_sync_blk;
    wire [18:0] proc_5_output_sync_blk;
    wire [18:0] proc_dep_vld_vec_5;
    reg [18:0] proc_dep_vld_vec_5_reg;
    wire [18:0] in_chan_dep_vld_vec_5;
    wire [664:0] in_chan_dep_data_vec_5;
    wire [18:0] token_in_vec_5;
    wire [18:0] out_chan_dep_vld_vec_5;
    wire [34:0] out_chan_dep_data_5;
    wire [18:0] token_out_vec_5;
    wire dl_detect_out_5;
    wire dep_chan_vld_0_5;
    wire [34:0] dep_chan_data_0_5;
    wire token_0_5;
    wire dep_chan_vld_1_5;
    wire [34:0] dep_chan_data_1_5;
    wire token_1_5;
    wire dep_chan_vld_2_5;
    wire [34:0] dep_chan_data_2_5;
    wire token_2_5;
    wire dep_chan_vld_3_5;
    wire [34:0] dep_chan_data_3_5;
    wire token_3_5;
    wire dep_chan_vld_4_5;
    wire [34:0] dep_chan_data_4_5;
    wire token_4_5;
    wire dep_chan_vld_6_5;
    wire [34:0] dep_chan_data_6_5;
    wire token_6_5;
    wire dep_chan_vld_7_5;
    wire [34:0] dep_chan_data_7_5;
    wire token_7_5;
    wire dep_chan_vld_8_5;
    wire [34:0] dep_chan_data_8_5;
    wire token_8_5;
    wire dep_chan_vld_9_5;
    wire [34:0] dep_chan_data_9_5;
    wire token_9_5;
    wire dep_chan_vld_10_5;
    wire [34:0] dep_chan_data_10_5;
    wire token_10_5;
    wire dep_chan_vld_11_5;
    wire [34:0] dep_chan_data_11_5;
    wire token_11_5;
    wire dep_chan_vld_12_5;
    wire [34:0] dep_chan_data_12_5;
    wire token_12_5;
    wire dep_chan_vld_13_5;
    wire [34:0] dep_chan_data_13_5;
    wire token_13_5;
    wire dep_chan_vld_14_5;
    wire [34:0] dep_chan_data_14_5;
    wire token_14_5;
    wire dep_chan_vld_15_5;
    wire [34:0] dep_chan_data_15_5;
    wire token_15_5;
    wire dep_chan_vld_16_5;
    wire [34:0] dep_chan_data_16_5;
    wire token_16_5;
    wire dep_chan_vld_17_5;
    wire [34:0] dep_chan_data_17_5;
    wire token_17_5;
    wire dep_chan_vld_18_5;
    wire [34:0] dep_chan_data_18_5;
    wire token_18_5;
    wire dep_chan_vld_21_5;
    wire [34:0] dep_chan_data_21_5;
    wire token_21_5;
    wire [18:0] proc_6_data_FIFO_blk;
    wire [18:0] proc_6_data_PIPO_blk;
    wire [18:0] proc_6_start_FIFO_blk;
    wire [18:0] proc_6_TLF_FIFO_blk;
    wire [18:0] proc_6_input_sync_blk;
    wire [18:0] proc_6_output_sync_blk;
    wire [18:0] proc_dep_vld_vec_6;
    reg [18:0] proc_dep_vld_vec_6_reg;
    wire [18:0] in_chan_dep_vld_vec_6;
    wire [664:0] in_chan_dep_data_vec_6;
    wire [18:0] token_in_vec_6;
    wire [18:0] out_chan_dep_vld_vec_6;
    wire [34:0] out_chan_dep_data_6;
    wire [18:0] token_out_vec_6;
    wire dl_detect_out_6;
    wire dep_chan_vld_0_6;
    wire [34:0] dep_chan_data_0_6;
    wire token_0_6;
    wire dep_chan_vld_1_6;
    wire [34:0] dep_chan_data_1_6;
    wire token_1_6;
    wire dep_chan_vld_2_6;
    wire [34:0] dep_chan_data_2_6;
    wire token_2_6;
    wire dep_chan_vld_3_6;
    wire [34:0] dep_chan_data_3_6;
    wire token_3_6;
    wire dep_chan_vld_4_6;
    wire [34:0] dep_chan_data_4_6;
    wire token_4_6;
    wire dep_chan_vld_5_6;
    wire [34:0] dep_chan_data_5_6;
    wire token_5_6;
    wire dep_chan_vld_7_6;
    wire [34:0] dep_chan_data_7_6;
    wire token_7_6;
    wire dep_chan_vld_8_6;
    wire [34:0] dep_chan_data_8_6;
    wire token_8_6;
    wire dep_chan_vld_9_6;
    wire [34:0] dep_chan_data_9_6;
    wire token_9_6;
    wire dep_chan_vld_10_6;
    wire [34:0] dep_chan_data_10_6;
    wire token_10_6;
    wire dep_chan_vld_11_6;
    wire [34:0] dep_chan_data_11_6;
    wire token_11_6;
    wire dep_chan_vld_12_6;
    wire [34:0] dep_chan_data_12_6;
    wire token_12_6;
    wire dep_chan_vld_13_6;
    wire [34:0] dep_chan_data_13_6;
    wire token_13_6;
    wire dep_chan_vld_14_6;
    wire [34:0] dep_chan_data_14_6;
    wire token_14_6;
    wire dep_chan_vld_15_6;
    wire [34:0] dep_chan_data_15_6;
    wire token_15_6;
    wire dep_chan_vld_16_6;
    wire [34:0] dep_chan_data_16_6;
    wire token_16_6;
    wire dep_chan_vld_17_6;
    wire [34:0] dep_chan_data_17_6;
    wire token_17_6;
    wire dep_chan_vld_18_6;
    wire [34:0] dep_chan_data_18_6;
    wire token_18_6;
    wire dep_chan_vld_22_6;
    wire [34:0] dep_chan_data_22_6;
    wire token_22_6;
    wire [18:0] proc_7_data_FIFO_blk;
    wire [18:0] proc_7_data_PIPO_blk;
    wire [18:0] proc_7_start_FIFO_blk;
    wire [18:0] proc_7_TLF_FIFO_blk;
    wire [18:0] proc_7_input_sync_blk;
    wire [18:0] proc_7_output_sync_blk;
    wire [18:0] proc_dep_vld_vec_7;
    reg [18:0] proc_dep_vld_vec_7_reg;
    wire [18:0] in_chan_dep_vld_vec_7;
    wire [664:0] in_chan_dep_data_vec_7;
    wire [18:0] token_in_vec_7;
    wire [18:0] out_chan_dep_vld_vec_7;
    wire [34:0] out_chan_dep_data_7;
    wire [18:0] token_out_vec_7;
    wire dl_detect_out_7;
    wire dep_chan_vld_0_7;
    wire [34:0] dep_chan_data_0_7;
    wire token_0_7;
    wire dep_chan_vld_1_7;
    wire [34:0] dep_chan_data_1_7;
    wire token_1_7;
    wire dep_chan_vld_2_7;
    wire [34:0] dep_chan_data_2_7;
    wire token_2_7;
    wire dep_chan_vld_3_7;
    wire [34:0] dep_chan_data_3_7;
    wire token_3_7;
    wire dep_chan_vld_4_7;
    wire [34:0] dep_chan_data_4_7;
    wire token_4_7;
    wire dep_chan_vld_5_7;
    wire [34:0] dep_chan_data_5_7;
    wire token_5_7;
    wire dep_chan_vld_6_7;
    wire [34:0] dep_chan_data_6_7;
    wire token_6_7;
    wire dep_chan_vld_8_7;
    wire [34:0] dep_chan_data_8_7;
    wire token_8_7;
    wire dep_chan_vld_9_7;
    wire [34:0] dep_chan_data_9_7;
    wire token_9_7;
    wire dep_chan_vld_10_7;
    wire [34:0] dep_chan_data_10_7;
    wire token_10_7;
    wire dep_chan_vld_11_7;
    wire [34:0] dep_chan_data_11_7;
    wire token_11_7;
    wire dep_chan_vld_12_7;
    wire [34:0] dep_chan_data_12_7;
    wire token_12_7;
    wire dep_chan_vld_13_7;
    wire [34:0] dep_chan_data_13_7;
    wire token_13_7;
    wire dep_chan_vld_14_7;
    wire [34:0] dep_chan_data_14_7;
    wire token_14_7;
    wire dep_chan_vld_15_7;
    wire [34:0] dep_chan_data_15_7;
    wire token_15_7;
    wire dep_chan_vld_16_7;
    wire [34:0] dep_chan_data_16_7;
    wire token_16_7;
    wire dep_chan_vld_17_7;
    wire [34:0] dep_chan_data_17_7;
    wire token_17_7;
    wire dep_chan_vld_18_7;
    wire [34:0] dep_chan_data_18_7;
    wire token_18_7;
    wire dep_chan_vld_23_7;
    wire [34:0] dep_chan_data_23_7;
    wire token_23_7;
    wire [18:0] proc_8_data_FIFO_blk;
    wire [18:0] proc_8_data_PIPO_blk;
    wire [18:0] proc_8_start_FIFO_blk;
    wire [18:0] proc_8_TLF_FIFO_blk;
    wire [18:0] proc_8_input_sync_blk;
    wire [18:0] proc_8_output_sync_blk;
    wire [18:0] proc_dep_vld_vec_8;
    reg [18:0] proc_dep_vld_vec_8_reg;
    wire [18:0] in_chan_dep_vld_vec_8;
    wire [664:0] in_chan_dep_data_vec_8;
    wire [18:0] token_in_vec_8;
    wire [18:0] out_chan_dep_vld_vec_8;
    wire [34:0] out_chan_dep_data_8;
    wire [18:0] token_out_vec_8;
    wire dl_detect_out_8;
    wire dep_chan_vld_0_8;
    wire [34:0] dep_chan_data_0_8;
    wire token_0_8;
    wire dep_chan_vld_1_8;
    wire [34:0] dep_chan_data_1_8;
    wire token_1_8;
    wire dep_chan_vld_2_8;
    wire [34:0] dep_chan_data_2_8;
    wire token_2_8;
    wire dep_chan_vld_3_8;
    wire [34:0] dep_chan_data_3_8;
    wire token_3_8;
    wire dep_chan_vld_4_8;
    wire [34:0] dep_chan_data_4_8;
    wire token_4_8;
    wire dep_chan_vld_5_8;
    wire [34:0] dep_chan_data_5_8;
    wire token_5_8;
    wire dep_chan_vld_6_8;
    wire [34:0] dep_chan_data_6_8;
    wire token_6_8;
    wire dep_chan_vld_7_8;
    wire [34:0] dep_chan_data_7_8;
    wire token_7_8;
    wire dep_chan_vld_9_8;
    wire [34:0] dep_chan_data_9_8;
    wire token_9_8;
    wire dep_chan_vld_10_8;
    wire [34:0] dep_chan_data_10_8;
    wire token_10_8;
    wire dep_chan_vld_11_8;
    wire [34:0] dep_chan_data_11_8;
    wire token_11_8;
    wire dep_chan_vld_12_8;
    wire [34:0] dep_chan_data_12_8;
    wire token_12_8;
    wire dep_chan_vld_13_8;
    wire [34:0] dep_chan_data_13_8;
    wire token_13_8;
    wire dep_chan_vld_14_8;
    wire [34:0] dep_chan_data_14_8;
    wire token_14_8;
    wire dep_chan_vld_15_8;
    wire [34:0] dep_chan_data_15_8;
    wire token_15_8;
    wire dep_chan_vld_16_8;
    wire [34:0] dep_chan_data_16_8;
    wire token_16_8;
    wire dep_chan_vld_17_8;
    wire [34:0] dep_chan_data_17_8;
    wire token_17_8;
    wire dep_chan_vld_18_8;
    wire [34:0] dep_chan_data_18_8;
    wire token_18_8;
    wire dep_chan_vld_24_8;
    wire [34:0] dep_chan_data_24_8;
    wire token_24_8;
    wire [18:0] proc_9_data_FIFO_blk;
    wire [18:0] proc_9_data_PIPO_blk;
    wire [18:0] proc_9_start_FIFO_blk;
    wire [18:0] proc_9_TLF_FIFO_blk;
    wire [18:0] proc_9_input_sync_blk;
    wire [18:0] proc_9_output_sync_blk;
    wire [18:0] proc_dep_vld_vec_9;
    reg [18:0] proc_dep_vld_vec_9_reg;
    wire [18:0] in_chan_dep_vld_vec_9;
    wire [664:0] in_chan_dep_data_vec_9;
    wire [18:0] token_in_vec_9;
    wire [18:0] out_chan_dep_vld_vec_9;
    wire [34:0] out_chan_dep_data_9;
    wire [18:0] token_out_vec_9;
    wire dl_detect_out_9;
    wire dep_chan_vld_0_9;
    wire [34:0] dep_chan_data_0_9;
    wire token_0_9;
    wire dep_chan_vld_1_9;
    wire [34:0] dep_chan_data_1_9;
    wire token_1_9;
    wire dep_chan_vld_2_9;
    wire [34:0] dep_chan_data_2_9;
    wire token_2_9;
    wire dep_chan_vld_3_9;
    wire [34:0] dep_chan_data_3_9;
    wire token_3_9;
    wire dep_chan_vld_4_9;
    wire [34:0] dep_chan_data_4_9;
    wire token_4_9;
    wire dep_chan_vld_5_9;
    wire [34:0] dep_chan_data_5_9;
    wire token_5_9;
    wire dep_chan_vld_6_9;
    wire [34:0] dep_chan_data_6_9;
    wire token_6_9;
    wire dep_chan_vld_7_9;
    wire [34:0] dep_chan_data_7_9;
    wire token_7_9;
    wire dep_chan_vld_8_9;
    wire [34:0] dep_chan_data_8_9;
    wire token_8_9;
    wire dep_chan_vld_10_9;
    wire [34:0] dep_chan_data_10_9;
    wire token_10_9;
    wire dep_chan_vld_11_9;
    wire [34:0] dep_chan_data_11_9;
    wire token_11_9;
    wire dep_chan_vld_12_9;
    wire [34:0] dep_chan_data_12_9;
    wire token_12_9;
    wire dep_chan_vld_13_9;
    wire [34:0] dep_chan_data_13_9;
    wire token_13_9;
    wire dep_chan_vld_14_9;
    wire [34:0] dep_chan_data_14_9;
    wire token_14_9;
    wire dep_chan_vld_15_9;
    wire [34:0] dep_chan_data_15_9;
    wire token_15_9;
    wire dep_chan_vld_16_9;
    wire [34:0] dep_chan_data_16_9;
    wire token_16_9;
    wire dep_chan_vld_17_9;
    wire [34:0] dep_chan_data_17_9;
    wire token_17_9;
    wire dep_chan_vld_18_9;
    wire [34:0] dep_chan_data_18_9;
    wire token_18_9;
    wire dep_chan_vld_25_9;
    wire [34:0] dep_chan_data_25_9;
    wire token_25_9;
    wire [18:0] proc_10_data_FIFO_blk;
    wire [18:0] proc_10_data_PIPO_blk;
    wire [18:0] proc_10_start_FIFO_blk;
    wire [18:0] proc_10_TLF_FIFO_blk;
    wire [18:0] proc_10_input_sync_blk;
    wire [18:0] proc_10_output_sync_blk;
    wire [18:0] proc_dep_vld_vec_10;
    reg [18:0] proc_dep_vld_vec_10_reg;
    wire [18:0] in_chan_dep_vld_vec_10;
    wire [664:0] in_chan_dep_data_vec_10;
    wire [18:0] token_in_vec_10;
    wire [18:0] out_chan_dep_vld_vec_10;
    wire [34:0] out_chan_dep_data_10;
    wire [18:0] token_out_vec_10;
    wire dl_detect_out_10;
    wire dep_chan_vld_0_10;
    wire [34:0] dep_chan_data_0_10;
    wire token_0_10;
    wire dep_chan_vld_1_10;
    wire [34:0] dep_chan_data_1_10;
    wire token_1_10;
    wire dep_chan_vld_2_10;
    wire [34:0] dep_chan_data_2_10;
    wire token_2_10;
    wire dep_chan_vld_3_10;
    wire [34:0] dep_chan_data_3_10;
    wire token_3_10;
    wire dep_chan_vld_4_10;
    wire [34:0] dep_chan_data_4_10;
    wire token_4_10;
    wire dep_chan_vld_5_10;
    wire [34:0] dep_chan_data_5_10;
    wire token_5_10;
    wire dep_chan_vld_6_10;
    wire [34:0] dep_chan_data_6_10;
    wire token_6_10;
    wire dep_chan_vld_7_10;
    wire [34:0] dep_chan_data_7_10;
    wire token_7_10;
    wire dep_chan_vld_8_10;
    wire [34:0] dep_chan_data_8_10;
    wire token_8_10;
    wire dep_chan_vld_9_10;
    wire [34:0] dep_chan_data_9_10;
    wire token_9_10;
    wire dep_chan_vld_11_10;
    wire [34:0] dep_chan_data_11_10;
    wire token_11_10;
    wire dep_chan_vld_12_10;
    wire [34:0] dep_chan_data_12_10;
    wire token_12_10;
    wire dep_chan_vld_13_10;
    wire [34:0] dep_chan_data_13_10;
    wire token_13_10;
    wire dep_chan_vld_14_10;
    wire [34:0] dep_chan_data_14_10;
    wire token_14_10;
    wire dep_chan_vld_15_10;
    wire [34:0] dep_chan_data_15_10;
    wire token_15_10;
    wire dep_chan_vld_16_10;
    wire [34:0] dep_chan_data_16_10;
    wire token_16_10;
    wire dep_chan_vld_17_10;
    wire [34:0] dep_chan_data_17_10;
    wire token_17_10;
    wire dep_chan_vld_18_10;
    wire [34:0] dep_chan_data_18_10;
    wire token_18_10;
    wire dep_chan_vld_26_10;
    wire [34:0] dep_chan_data_26_10;
    wire token_26_10;
    wire [18:0] proc_11_data_FIFO_blk;
    wire [18:0] proc_11_data_PIPO_blk;
    wire [18:0] proc_11_start_FIFO_blk;
    wire [18:0] proc_11_TLF_FIFO_blk;
    wire [18:0] proc_11_input_sync_blk;
    wire [18:0] proc_11_output_sync_blk;
    wire [18:0] proc_dep_vld_vec_11;
    reg [18:0] proc_dep_vld_vec_11_reg;
    wire [18:0] in_chan_dep_vld_vec_11;
    wire [664:0] in_chan_dep_data_vec_11;
    wire [18:0] token_in_vec_11;
    wire [18:0] out_chan_dep_vld_vec_11;
    wire [34:0] out_chan_dep_data_11;
    wire [18:0] token_out_vec_11;
    wire dl_detect_out_11;
    wire dep_chan_vld_0_11;
    wire [34:0] dep_chan_data_0_11;
    wire token_0_11;
    wire dep_chan_vld_1_11;
    wire [34:0] dep_chan_data_1_11;
    wire token_1_11;
    wire dep_chan_vld_2_11;
    wire [34:0] dep_chan_data_2_11;
    wire token_2_11;
    wire dep_chan_vld_3_11;
    wire [34:0] dep_chan_data_3_11;
    wire token_3_11;
    wire dep_chan_vld_4_11;
    wire [34:0] dep_chan_data_4_11;
    wire token_4_11;
    wire dep_chan_vld_5_11;
    wire [34:0] dep_chan_data_5_11;
    wire token_5_11;
    wire dep_chan_vld_6_11;
    wire [34:0] dep_chan_data_6_11;
    wire token_6_11;
    wire dep_chan_vld_7_11;
    wire [34:0] dep_chan_data_7_11;
    wire token_7_11;
    wire dep_chan_vld_8_11;
    wire [34:0] dep_chan_data_8_11;
    wire token_8_11;
    wire dep_chan_vld_9_11;
    wire [34:0] dep_chan_data_9_11;
    wire token_9_11;
    wire dep_chan_vld_10_11;
    wire [34:0] dep_chan_data_10_11;
    wire token_10_11;
    wire dep_chan_vld_12_11;
    wire [34:0] dep_chan_data_12_11;
    wire token_12_11;
    wire dep_chan_vld_13_11;
    wire [34:0] dep_chan_data_13_11;
    wire token_13_11;
    wire dep_chan_vld_14_11;
    wire [34:0] dep_chan_data_14_11;
    wire token_14_11;
    wire dep_chan_vld_15_11;
    wire [34:0] dep_chan_data_15_11;
    wire token_15_11;
    wire dep_chan_vld_16_11;
    wire [34:0] dep_chan_data_16_11;
    wire token_16_11;
    wire dep_chan_vld_17_11;
    wire [34:0] dep_chan_data_17_11;
    wire token_17_11;
    wire dep_chan_vld_18_11;
    wire [34:0] dep_chan_data_18_11;
    wire token_18_11;
    wire dep_chan_vld_27_11;
    wire [34:0] dep_chan_data_27_11;
    wire token_27_11;
    wire [18:0] proc_12_data_FIFO_blk;
    wire [18:0] proc_12_data_PIPO_blk;
    wire [18:0] proc_12_start_FIFO_blk;
    wire [18:0] proc_12_TLF_FIFO_blk;
    wire [18:0] proc_12_input_sync_blk;
    wire [18:0] proc_12_output_sync_blk;
    wire [18:0] proc_dep_vld_vec_12;
    reg [18:0] proc_dep_vld_vec_12_reg;
    wire [18:0] in_chan_dep_vld_vec_12;
    wire [664:0] in_chan_dep_data_vec_12;
    wire [18:0] token_in_vec_12;
    wire [18:0] out_chan_dep_vld_vec_12;
    wire [34:0] out_chan_dep_data_12;
    wire [18:0] token_out_vec_12;
    wire dl_detect_out_12;
    wire dep_chan_vld_0_12;
    wire [34:0] dep_chan_data_0_12;
    wire token_0_12;
    wire dep_chan_vld_1_12;
    wire [34:0] dep_chan_data_1_12;
    wire token_1_12;
    wire dep_chan_vld_2_12;
    wire [34:0] dep_chan_data_2_12;
    wire token_2_12;
    wire dep_chan_vld_3_12;
    wire [34:0] dep_chan_data_3_12;
    wire token_3_12;
    wire dep_chan_vld_4_12;
    wire [34:0] dep_chan_data_4_12;
    wire token_4_12;
    wire dep_chan_vld_5_12;
    wire [34:0] dep_chan_data_5_12;
    wire token_5_12;
    wire dep_chan_vld_6_12;
    wire [34:0] dep_chan_data_6_12;
    wire token_6_12;
    wire dep_chan_vld_7_12;
    wire [34:0] dep_chan_data_7_12;
    wire token_7_12;
    wire dep_chan_vld_8_12;
    wire [34:0] dep_chan_data_8_12;
    wire token_8_12;
    wire dep_chan_vld_9_12;
    wire [34:0] dep_chan_data_9_12;
    wire token_9_12;
    wire dep_chan_vld_10_12;
    wire [34:0] dep_chan_data_10_12;
    wire token_10_12;
    wire dep_chan_vld_11_12;
    wire [34:0] dep_chan_data_11_12;
    wire token_11_12;
    wire dep_chan_vld_13_12;
    wire [34:0] dep_chan_data_13_12;
    wire token_13_12;
    wire dep_chan_vld_14_12;
    wire [34:0] dep_chan_data_14_12;
    wire token_14_12;
    wire dep_chan_vld_15_12;
    wire [34:0] dep_chan_data_15_12;
    wire token_15_12;
    wire dep_chan_vld_16_12;
    wire [34:0] dep_chan_data_16_12;
    wire token_16_12;
    wire dep_chan_vld_17_12;
    wire [34:0] dep_chan_data_17_12;
    wire token_17_12;
    wire dep_chan_vld_18_12;
    wire [34:0] dep_chan_data_18_12;
    wire token_18_12;
    wire dep_chan_vld_28_12;
    wire [34:0] dep_chan_data_28_12;
    wire token_28_12;
    wire [18:0] proc_13_data_FIFO_blk;
    wire [18:0] proc_13_data_PIPO_blk;
    wire [18:0] proc_13_start_FIFO_blk;
    wire [18:0] proc_13_TLF_FIFO_blk;
    wire [18:0] proc_13_input_sync_blk;
    wire [18:0] proc_13_output_sync_blk;
    wire [18:0] proc_dep_vld_vec_13;
    reg [18:0] proc_dep_vld_vec_13_reg;
    wire [18:0] in_chan_dep_vld_vec_13;
    wire [664:0] in_chan_dep_data_vec_13;
    wire [18:0] token_in_vec_13;
    wire [18:0] out_chan_dep_vld_vec_13;
    wire [34:0] out_chan_dep_data_13;
    wire [18:0] token_out_vec_13;
    wire dl_detect_out_13;
    wire dep_chan_vld_0_13;
    wire [34:0] dep_chan_data_0_13;
    wire token_0_13;
    wire dep_chan_vld_1_13;
    wire [34:0] dep_chan_data_1_13;
    wire token_1_13;
    wire dep_chan_vld_2_13;
    wire [34:0] dep_chan_data_2_13;
    wire token_2_13;
    wire dep_chan_vld_3_13;
    wire [34:0] dep_chan_data_3_13;
    wire token_3_13;
    wire dep_chan_vld_4_13;
    wire [34:0] dep_chan_data_4_13;
    wire token_4_13;
    wire dep_chan_vld_5_13;
    wire [34:0] dep_chan_data_5_13;
    wire token_5_13;
    wire dep_chan_vld_6_13;
    wire [34:0] dep_chan_data_6_13;
    wire token_6_13;
    wire dep_chan_vld_7_13;
    wire [34:0] dep_chan_data_7_13;
    wire token_7_13;
    wire dep_chan_vld_8_13;
    wire [34:0] dep_chan_data_8_13;
    wire token_8_13;
    wire dep_chan_vld_9_13;
    wire [34:0] dep_chan_data_9_13;
    wire token_9_13;
    wire dep_chan_vld_10_13;
    wire [34:0] dep_chan_data_10_13;
    wire token_10_13;
    wire dep_chan_vld_11_13;
    wire [34:0] dep_chan_data_11_13;
    wire token_11_13;
    wire dep_chan_vld_12_13;
    wire [34:0] dep_chan_data_12_13;
    wire token_12_13;
    wire dep_chan_vld_14_13;
    wire [34:0] dep_chan_data_14_13;
    wire token_14_13;
    wire dep_chan_vld_15_13;
    wire [34:0] dep_chan_data_15_13;
    wire token_15_13;
    wire dep_chan_vld_16_13;
    wire [34:0] dep_chan_data_16_13;
    wire token_16_13;
    wire dep_chan_vld_17_13;
    wire [34:0] dep_chan_data_17_13;
    wire token_17_13;
    wire dep_chan_vld_18_13;
    wire [34:0] dep_chan_data_18_13;
    wire token_18_13;
    wire dep_chan_vld_29_13;
    wire [34:0] dep_chan_data_29_13;
    wire token_29_13;
    wire [18:0] proc_14_data_FIFO_blk;
    wire [18:0] proc_14_data_PIPO_blk;
    wire [18:0] proc_14_start_FIFO_blk;
    wire [18:0] proc_14_TLF_FIFO_blk;
    wire [18:0] proc_14_input_sync_blk;
    wire [18:0] proc_14_output_sync_blk;
    wire [18:0] proc_dep_vld_vec_14;
    reg [18:0] proc_dep_vld_vec_14_reg;
    wire [18:0] in_chan_dep_vld_vec_14;
    wire [664:0] in_chan_dep_data_vec_14;
    wire [18:0] token_in_vec_14;
    wire [18:0] out_chan_dep_vld_vec_14;
    wire [34:0] out_chan_dep_data_14;
    wire [18:0] token_out_vec_14;
    wire dl_detect_out_14;
    wire dep_chan_vld_0_14;
    wire [34:0] dep_chan_data_0_14;
    wire token_0_14;
    wire dep_chan_vld_1_14;
    wire [34:0] dep_chan_data_1_14;
    wire token_1_14;
    wire dep_chan_vld_2_14;
    wire [34:0] dep_chan_data_2_14;
    wire token_2_14;
    wire dep_chan_vld_3_14;
    wire [34:0] dep_chan_data_3_14;
    wire token_3_14;
    wire dep_chan_vld_4_14;
    wire [34:0] dep_chan_data_4_14;
    wire token_4_14;
    wire dep_chan_vld_5_14;
    wire [34:0] dep_chan_data_5_14;
    wire token_5_14;
    wire dep_chan_vld_6_14;
    wire [34:0] dep_chan_data_6_14;
    wire token_6_14;
    wire dep_chan_vld_7_14;
    wire [34:0] dep_chan_data_7_14;
    wire token_7_14;
    wire dep_chan_vld_8_14;
    wire [34:0] dep_chan_data_8_14;
    wire token_8_14;
    wire dep_chan_vld_9_14;
    wire [34:0] dep_chan_data_9_14;
    wire token_9_14;
    wire dep_chan_vld_10_14;
    wire [34:0] dep_chan_data_10_14;
    wire token_10_14;
    wire dep_chan_vld_11_14;
    wire [34:0] dep_chan_data_11_14;
    wire token_11_14;
    wire dep_chan_vld_12_14;
    wire [34:0] dep_chan_data_12_14;
    wire token_12_14;
    wire dep_chan_vld_13_14;
    wire [34:0] dep_chan_data_13_14;
    wire token_13_14;
    wire dep_chan_vld_15_14;
    wire [34:0] dep_chan_data_15_14;
    wire token_15_14;
    wire dep_chan_vld_16_14;
    wire [34:0] dep_chan_data_16_14;
    wire token_16_14;
    wire dep_chan_vld_17_14;
    wire [34:0] dep_chan_data_17_14;
    wire token_17_14;
    wire dep_chan_vld_18_14;
    wire [34:0] dep_chan_data_18_14;
    wire token_18_14;
    wire dep_chan_vld_30_14;
    wire [34:0] dep_chan_data_30_14;
    wire token_30_14;
    wire [18:0] proc_15_data_FIFO_blk;
    wire [18:0] proc_15_data_PIPO_blk;
    wire [18:0] proc_15_start_FIFO_blk;
    wire [18:0] proc_15_TLF_FIFO_blk;
    wire [18:0] proc_15_input_sync_blk;
    wire [18:0] proc_15_output_sync_blk;
    wire [18:0] proc_dep_vld_vec_15;
    reg [18:0] proc_dep_vld_vec_15_reg;
    wire [18:0] in_chan_dep_vld_vec_15;
    wire [664:0] in_chan_dep_data_vec_15;
    wire [18:0] token_in_vec_15;
    wire [18:0] out_chan_dep_vld_vec_15;
    wire [34:0] out_chan_dep_data_15;
    wire [18:0] token_out_vec_15;
    wire dl_detect_out_15;
    wire dep_chan_vld_0_15;
    wire [34:0] dep_chan_data_0_15;
    wire token_0_15;
    wire dep_chan_vld_1_15;
    wire [34:0] dep_chan_data_1_15;
    wire token_1_15;
    wire dep_chan_vld_2_15;
    wire [34:0] dep_chan_data_2_15;
    wire token_2_15;
    wire dep_chan_vld_3_15;
    wire [34:0] dep_chan_data_3_15;
    wire token_3_15;
    wire dep_chan_vld_4_15;
    wire [34:0] dep_chan_data_4_15;
    wire token_4_15;
    wire dep_chan_vld_5_15;
    wire [34:0] dep_chan_data_5_15;
    wire token_5_15;
    wire dep_chan_vld_6_15;
    wire [34:0] dep_chan_data_6_15;
    wire token_6_15;
    wire dep_chan_vld_7_15;
    wire [34:0] dep_chan_data_7_15;
    wire token_7_15;
    wire dep_chan_vld_8_15;
    wire [34:0] dep_chan_data_8_15;
    wire token_8_15;
    wire dep_chan_vld_9_15;
    wire [34:0] dep_chan_data_9_15;
    wire token_9_15;
    wire dep_chan_vld_10_15;
    wire [34:0] dep_chan_data_10_15;
    wire token_10_15;
    wire dep_chan_vld_11_15;
    wire [34:0] dep_chan_data_11_15;
    wire token_11_15;
    wire dep_chan_vld_12_15;
    wire [34:0] dep_chan_data_12_15;
    wire token_12_15;
    wire dep_chan_vld_13_15;
    wire [34:0] dep_chan_data_13_15;
    wire token_13_15;
    wire dep_chan_vld_14_15;
    wire [34:0] dep_chan_data_14_15;
    wire token_14_15;
    wire dep_chan_vld_16_15;
    wire [34:0] dep_chan_data_16_15;
    wire token_16_15;
    wire dep_chan_vld_17_15;
    wire [34:0] dep_chan_data_17_15;
    wire token_17_15;
    wire dep_chan_vld_18_15;
    wire [34:0] dep_chan_data_18_15;
    wire token_18_15;
    wire dep_chan_vld_31_15;
    wire [34:0] dep_chan_data_31_15;
    wire token_31_15;
    wire [18:0] proc_16_data_FIFO_blk;
    wire [18:0] proc_16_data_PIPO_blk;
    wire [18:0] proc_16_start_FIFO_blk;
    wire [18:0] proc_16_TLF_FIFO_blk;
    wire [18:0] proc_16_input_sync_blk;
    wire [18:0] proc_16_output_sync_blk;
    wire [18:0] proc_dep_vld_vec_16;
    reg [18:0] proc_dep_vld_vec_16_reg;
    wire [18:0] in_chan_dep_vld_vec_16;
    wire [664:0] in_chan_dep_data_vec_16;
    wire [18:0] token_in_vec_16;
    wire [18:0] out_chan_dep_vld_vec_16;
    wire [34:0] out_chan_dep_data_16;
    wire [18:0] token_out_vec_16;
    wire dl_detect_out_16;
    wire dep_chan_vld_0_16;
    wire [34:0] dep_chan_data_0_16;
    wire token_0_16;
    wire dep_chan_vld_1_16;
    wire [34:0] dep_chan_data_1_16;
    wire token_1_16;
    wire dep_chan_vld_2_16;
    wire [34:0] dep_chan_data_2_16;
    wire token_2_16;
    wire dep_chan_vld_3_16;
    wire [34:0] dep_chan_data_3_16;
    wire token_3_16;
    wire dep_chan_vld_4_16;
    wire [34:0] dep_chan_data_4_16;
    wire token_4_16;
    wire dep_chan_vld_5_16;
    wire [34:0] dep_chan_data_5_16;
    wire token_5_16;
    wire dep_chan_vld_6_16;
    wire [34:0] dep_chan_data_6_16;
    wire token_6_16;
    wire dep_chan_vld_7_16;
    wire [34:0] dep_chan_data_7_16;
    wire token_7_16;
    wire dep_chan_vld_8_16;
    wire [34:0] dep_chan_data_8_16;
    wire token_8_16;
    wire dep_chan_vld_9_16;
    wire [34:0] dep_chan_data_9_16;
    wire token_9_16;
    wire dep_chan_vld_10_16;
    wire [34:0] dep_chan_data_10_16;
    wire token_10_16;
    wire dep_chan_vld_11_16;
    wire [34:0] dep_chan_data_11_16;
    wire token_11_16;
    wire dep_chan_vld_12_16;
    wire [34:0] dep_chan_data_12_16;
    wire token_12_16;
    wire dep_chan_vld_13_16;
    wire [34:0] dep_chan_data_13_16;
    wire token_13_16;
    wire dep_chan_vld_14_16;
    wire [34:0] dep_chan_data_14_16;
    wire token_14_16;
    wire dep_chan_vld_15_16;
    wire [34:0] dep_chan_data_15_16;
    wire token_15_16;
    wire dep_chan_vld_17_16;
    wire [34:0] dep_chan_data_17_16;
    wire token_17_16;
    wire dep_chan_vld_18_16;
    wire [34:0] dep_chan_data_18_16;
    wire token_18_16;
    wire dep_chan_vld_32_16;
    wire [34:0] dep_chan_data_32_16;
    wire token_32_16;
    wire [18:0] proc_17_data_FIFO_blk;
    wire [18:0] proc_17_data_PIPO_blk;
    wire [18:0] proc_17_start_FIFO_blk;
    wire [18:0] proc_17_TLF_FIFO_blk;
    wire [18:0] proc_17_input_sync_blk;
    wire [18:0] proc_17_output_sync_blk;
    wire [18:0] proc_dep_vld_vec_17;
    reg [18:0] proc_dep_vld_vec_17_reg;
    wire [18:0] in_chan_dep_vld_vec_17;
    wire [664:0] in_chan_dep_data_vec_17;
    wire [18:0] token_in_vec_17;
    wire [18:0] out_chan_dep_vld_vec_17;
    wire [34:0] out_chan_dep_data_17;
    wire [18:0] token_out_vec_17;
    wire dl_detect_out_17;
    wire dep_chan_vld_0_17;
    wire [34:0] dep_chan_data_0_17;
    wire token_0_17;
    wire dep_chan_vld_1_17;
    wire [34:0] dep_chan_data_1_17;
    wire token_1_17;
    wire dep_chan_vld_2_17;
    wire [34:0] dep_chan_data_2_17;
    wire token_2_17;
    wire dep_chan_vld_3_17;
    wire [34:0] dep_chan_data_3_17;
    wire token_3_17;
    wire dep_chan_vld_4_17;
    wire [34:0] dep_chan_data_4_17;
    wire token_4_17;
    wire dep_chan_vld_5_17;
    wire [34:0] dep_chan_data_5_17;
    wire token_5_17;
    wire dep_chan_vld_6_17;
    wire [34:0] dep_chan_data_6_17;
    wire token_6_17;
    wire dep_chan_vld_7_17;
    wire [34:0] dep_chan_data_7_17;
    wire token_7_17;
    wire dep_chan_vld_8_17;
    wire [34:0] dep_chan_data_8_17;
    wire token_8_17;
    wire dep_chan_vld_9_17;
    wire [34:0] dep_chan_data_9_17;
    wire token_9_17;
    wire dep_chan_vld_10_17;
    wire [34:0] dep_chan_data_10_17;
    wire token_10_17;
    wire dep_chan_vld_11_17;
    wire [34:0] dep_chan_data_11_17;
    wire token_11_17;
    wire dep_chan_vld_12_17;
    wire [34:0] dep_chan_data_12_17;
    wire token_12_17;
    wire dep_chan_vld_13_17;
    wire [34:0] dep_chan_data_13_17;
    wire token_13_17;
    wire dep_chan_vld_14_17;
    wire [34:0] dep_chan_data_14_17;
    wire token_14_17;
    wire dep_chan_vld_15_17;
    wire [34:0] dep_chan_data_15_17;
    wire token_15_17;
    wire dep_chan_vld_16_17;
    wire [34:0] dep_chan_data_16_17;
    wire token_16_17;
    wire dep_chan_vld_18_17;
    wire [34:0] dep_chan_data_18_17;
    wire token_18_17;
    wire dep_chan_vld_33_17;
    wire [34:0] dep_chan_data_33_17;
    wire token_33_17;
    wire [18:0] proc_18_data_FIFO_blk;
    wire [18:0] proc_18_data_PIPO_blk;
    wire [18:0] proc_18_start_FIFO_blk;
    wire [18:0] proc_18_TLF_FIFO_blk;
    wire [18:0] proc_18_input_sync_blk;
    wire [18:0] proc_18_output_sync_blk;
    wire [18:0] proc_dep_vld_vec_18;
    reg [18:0] proc_dep_vld_vec_18_reg;
    wire [18:0] in_chan_dep_vld_vec_18;
    wire [664:0] in_chan_dep_data_vec_18;
    wire [18:0] token_in_vec_18;
    wire [18:0] out_chan_dep_vld_vec_18;
    wire [34:0] out_chan_dep_data_18;
    wire [18:0] token_out_vec_18;
    wire dl_detect_out_18;
    wire dep_chan_vld_0_18;
    wire [34:0] dep_chan_data_0_18;
    wire token_0_18;
    wire dep_chan_vld_1_18;
    wire [34:0] dep_chan_data_1_18;
    wire token_1_18;
    wire dep_chan_vld_2_18;
    wire [34:0] dep_chan_data_2_18;
    wire token_2_18;
    wire dep_chan_vld_3_18;
    wire [34:0] dep_chan_data_3_18;
    wire token_3_18;
    wire dep_chan_vld_4_18;
    wire [34:0] dep_chan_data_4_18;
    wire token_4_18;
    wire dep_chan_vld_5_18;
    wire [34:0] dep_chan_data_5_18;
    wire token_5_18;
    wire dep_chan_vld_6_18;
    wire [34:0] dep_chan_data_6_18;
    wire token_6_18;
    wire dep_chan_vld_7_18;
    wire [34:0] dep_chan_data_7_18;
    wire token_7_18;
    wire dep_chan_vld_8_18;
    wire [34:0] dep_chan_data_8_18;
    wire token_8_18;
    wire dep_chan_vld_9_18;
    wire [34:0] dep_chan_data_9_18;
    wire token_9_18;
    wire dep_chan_vld_10_18;
    wire [34:0] dep_chan_data_10_18;
    wire token_10_18;
    wire dep_chan_vld_11_18;
    wire [34:0] dep_chan_data_11_18;
    wire token_11_18;
    wire dep_chan_vld_12_18;
    wire [34:0] dep_chan_data_12_18;
    wire token_12_18;
    wire dep_chan_vld_13_18;
    wire [34:0] dep_chan_data_13_18;
    wire token_13_18;
    wire dep_chan_vld_14_18;
    wire [34:0] dep_chan_data_14_18;
    wire token_14_18;
    wire dep_chan_vld_15_18;
    wire [34:0] dep_chan_data_15_18;
    wire token_15_18;
    wire dep_chan_vld_16_18;
    wire [34:0] dep_chan_data_16_18;
    wire token_16_18;
    wire dep_chan_vld_17_18;
    wire [34:0] dep_chan_data_17_18;
    wire token_17_18;
    wire dep_chan_vld_34_18;
    wire [34:0] dep_chan_data_34_18;
    wire token_34_18;
    wire [16:0] proc_19_data_FIFO_blk;
    wire [16:0] proc_19_data_PIPO_blk;
    wire [16:0] proc_19_start_FIFO_blk;
    wire [16:0] proc_19_TLF_FIFO_blk;
    wire [16:0] proc_19_input_sync_blk;
    wire [16:0] proc_19_output_sync_blk;
    wire [16:0] proc_dep_vld_vec_19;
    reg [16:0] proc_dep_vld_vec_19_reg;
    wire [16:0] in_chan_dep_vld_vec_19;
    wire [594:0] in_chan_dep_data_vec_19;
    wire [16:0] token_in_vec_19;
    wire [16:0] out_chan_dep_vld_vec_19;
    wire [34:0] out_chan_dep_data_19;
    wire [16:0] token_out_vec_19;
    wire dl_detect_out_19;
    wire dep_chan_vld_0_19;
    wire [34:0] dep_chan_data_0_19;
    wire token_0_19;
    wire dep_chan_vld_3_19;
    wire [34:0] dep_chan_data_3_19;
    wire token_3_19;
    wire dep_chan_vld_20_19;
    wire [34:0] dep_chan_data_20_19;
    wire token_20_19;
    wire dep_chan_vld_21_19;
    wire [34:0] dep_chan_data_21_19;
    wire token_21_19;
    wire dep_chan_vld_22_19;
    wire [34:0] dep_chan_data_22_19;
    wire token_22_19;
    wire dep_chan_vld_23_19;
    wire [34:0] dep_chan_data_23_19;
    wire token_23_19;
    wire dep_chan_vld_24_19;
    wire [34:0] dep_chan_data_24_19;
    wire token_24_19;
    wire dep_chan_vld_25_19;
    wire [34:0] dep_chan_data_25_19;
    wire token_25_19;
    wire dep_chan_vld_26_19;
    wire [34:0] dep_chan_data_26_19;
    wire token_26_19;
    wire dep_chan_vld_27_19;
    wire [34:0] dep_chan_data_27_19;
    wire token_27_19;
    wire dep_chan_vld_28_19;
    wire [34:0] dep_chan_data_28_19;
    wire token_28_19;
    wire dep_chan_vld_29_19;
    wire [34:0] dep_chan_data_29_19;
    wire token_29_19;
    wire dep_chan_vld_30_19;
    wire [34:0] dep_chan_data_30_19;
    wire token_30_19;
    wire dep_chan_vld_31_19;
    wire [34:0] dep_chan_data_31_19;
    wire token_31_19;
    wire dep_chan_vld_32_19;
    wire [34:0] dep_chan_data_32_19;
    wire token_32_19;
    wire dep_chan_vld_33_19;
    wire [34:0] dep_chan_data_33_19;
    wire token_33_19;
    wire dep_chan_vld_34_19;
    wire [34:0] dep_chan_data_34_19;
    wire token_34_19;
    wire [16:0] proc_20_data_FIFO_blk;
    wire [16:0] proc_20_data_PIPO_blk;
    wire [16:0] proc_20_start_FIFO_blk;
    wire [16:0] proc_20_TLF_FIFO_blk;
    wire [16:0] proc_20_input_sync_blk;
    wire [16:0] proc_20_output_sync_blk;
    wire [16:0] proc_dep_vld_vec_20;
    reg [16:0] proc_dep_vld_vec_20_reg;
    wire [16:0] in_chan_dep_vld_vec_20;
    wire [594:0] in_chan_dep_data_vec_20;
    wire [16:0] token_in_vec_20;
    wire [16:0] out_chan_dep_vld_vec_20;
    wire [34:0] out_chan_dep_data_20;
    wire [16:0] token_out_vec_20;
    wire dl_detect_out_20;
    wire dep_chan_vld_0_20;
    wire [34:0] dep_chan_data_0_20;
    wire token_0_20;
    wire dep_chan_vld_4_20;
    wire [34:0] dep_chan_data_4_20;
    wire token_4_20;
    wire dep_chan_vld_19_20;
    wire [34:0] dep_chan_data_19_20;
    wire token_19_20;
    wire dep_chan_vld_21_20;
    wire [34:0] dep_chan_data_21_20;
    wire token_21_20;
    wire dep_chan_vld_22_20;
    wire [34:0] dep_chan_data_22_20;
    wire token_22_20;
    wire dep_chan_vld_23_20;
    wire [34:0] dep_chan_data_23_20;
    wire token_23_20;
    wire dep_chan_vld_24_20;
    wire [34:0] dep_chan_data_24_20;
    wire token_24_20;
    wire dep_chan_vld_25_20;
    wire [34:0] dep_chan_data_25_20;
    wire token_25_20;
    wire dep_chan_vld_26_20;
    wire [34:0] dep_chan_data_26_20;
    wire token_26_20;
    wire dep_chan_vld_27_20;
    wire [34:0] dep_chan_data_27_20;
    wire token_27_20;
    wire dep_chan_vld_28_20;
    wire [34:0] dep_chan_data_28_20;
    wire token_28_20;
    wire dep_chan_vld_29_20;
    wire [34:0] dep_chan_data_29_20;
    wire token_29_20;
    wire dep_chan_vld_30_20;
    wire [34:0] dep_chan_data_30_20;
    wire token_30_20;
    wire dep_chan_vld_31_20;
    wire [34:0] dep_chan_data_31_20;
    wire token_31_20;
    wire dep_chan_vld_32_20;
    wire [34:0] dep_chan_data_32_20;
    wire token_32_20;
    wire dep_chan_vld_33_20;
    wire [34:0] dep_chan_data_33_20;
    wire token_33_20;
    wire dep_chan_vld_34_20;
    wire [34:0] dep_chan_data_34_20;
    wire token_34_20;
    wire [16:0] proc_21_data_FIFO_blk;
    wire [16:0] proc_21_data_PIPO_blk;
    wire [16:0] proc_21_start_FIFO_blk;
    wire [16:0] proc_21_TLF_FIFO_blk;
    wire [16:0] proc_21_input_sync_blk;
    wire [16:0] proc_21_output_sync_blk;
    wire [16:0] proc_dep_vld_vec_21;
    reg [16:0] proc_dep_vld_vec_21_reg;
    wire [16:0] in_chan_dep_vld_vec_21;
    wire [594:0] in_chan_dep_data_vec_21;
    wire [16:0] token_in_vec_21;
    wire [16:0] out_chan_dep_vld_vec_21;
    wire [34:0] out_chan_dep_data_21;
    wire [16:0] token_out_vec_21;
    wire dl_detect_out_21;
    wire dep_chan_vld_0_21;
    wire [34:0] dep_chan_data_0_21;
    wire token_0_21;
    wire dep_chan_vld_5_21;
    wire [34:0] dep_chan_data_5_21;
    wire token_5_21;
    wire dep_chan_vld_19_21;
    wire [34:0] dep_chan_data_19_21;
    wire token_19_21;
    wire dep_chan_vld_20_21;
    wire [34:0] dep_chan_data_20_21;
    wire token_20_21;
    wire dep_chan_vld_22_21;
    wire [34:0] dep_chan_data_22_21;
    wire token_22_21;
    wire dep_chan_vld_23_21;
    wire [34:0] dep_chan_data_23_21;
    wire token_23_21;
    wire dep_chan_vld_24_21;
    wire [34:0] dep_chan_data_24_21;
    wire token_24_21;
    wire dep_chan_vld_25_21;
    wire [34:0] dep_chan_data_25_21;
    wire token_25_21;
    wire dep_chan_vld_26_21;
    wire [34:0] dep_chan_data_26_21;
    wire token_26_21;
    wire dep_chan_vld_27_21;
    wire [34:0] dep_chan_data_27_21;
    wire token_27_21;
    wire dep_chan_vld_28_21;
    wire [34:0] dep_chan_data_28_21;
    wire token_28_21;
    wire dep_chan_vld_29_21;
    wire [34:0] dep_chan_data_29_21;
    wire token_29_21;
    wire dep_chan_vld_30_21;
    wire [34:0] dep_chan_data_30_21;
    wire token_30_21;
    wire dep_chan_vld_31_21;
    wire [34:0] dep_chan_data_31_21;
    wire token_31_21;
    wire dep_chan_vld_32_21;
    wire [34:0] dep_chan_data_32_21;
    wire token_32_21;
    wire dep_chan_vld_33_21;
    wire [34:0] dep_chan_data_33_21;
    wire token_33_21;
    wire dep_chan_vld_34_21;
    wire [34:0] dep_chan_data_34_21;
    wire token_34_21;
    wire [16:0] proc_22_data_FIFO_blk;
    wire [16:0] proc_22_data_PIPO_blk;
    wire [16:0] proc_22_start_FIFO_blk;
    wire [16:0] proc_22_TLF_FIFO_blk;
    wire [16:0] proc_22_input_sync_blk;
    wire [16:0] proc_22_output_sync_blk;
    wire [16:0] proc_dep_vld_vec_22;
    reg [16:0] proc_dep_vld_vec_22_reg;
    wire [16:0] in_chan_dep_vld_vec_22;
    wire [594:0] in_chan_dep_data_vec_22;
    wire [16:0] token_in_vec_22;
    wire [16:0] out_chan_dep_vld_vec_22;
    wire [34:0] out_chan_dep_data_22;
    wire [16:0] token_out_vec_22;
    wire dl_detect_out_22;
    wire dep_chan_vld_0_22;
    wire [34:0] dep_chan_data_0_22;
    wire token_0_22;
    wire dep_chan_vld_6_22;
    wire [34:0] dep_chan_data_6_22;
    wire token_6_22;
    wire dep_chan_vld_19_22;
    wire [34:0] dep_chan_data_19_22;
    wire token_19_22;
    wire dep_chan_vld_20_22;
    wire [34:0] dep_chan_data_20_22;
    wire token_20_22;
    wire dep_chan_vld_21_22;
    wire [34:0] dep_chan_data_21_22;
    wire token_21_22;
    wire dep_chan_vld_23_22;
    wire [34:0] dep_chan_data_23_22;
    wire token_23_22;
    wire dep_chan_vld_24_22;
    wire [34:0] dep_chan_data_24_22;
    wire token_24_22;
    wire dep_chan_vld_25_22;
    wire [34:0] dep_chan_data_25_22;
    wire token_25_22;
    wire dep_chan_vld_26_22;
    wire [34:0] dep_chan_data_26_22;
    wire token_26_22;
    wire dep_chan_vld_27_22;
    wire [34:0] dep_chan_data_27_22;
    wire token_27_22;
    wire dep_chan_vld_28_22;
    wire [34:0] dep_chan_data_28_22;
    wire token_28_22;
    wire dep_chan_vld_29_22;
    wire [34:0] dep_chan_data_29_22;
    wire token_29_22;
    wire dep_chan_vld_30_22;
    wire [34:0] dep_chan_data_30_22;
    wire token_30_22;
    wire dep_chan_vld_31_22;
    wire [34:0] dep_chan_data_31_22;
    wire token_31_22;
    wire dep_chan_vld_32_22;
    wire [34:0] dep_chan_data_32_22;
    wire token_32_22;
    wire dep_chan_vld_33_22;
    wire [34:0] dep_chan_data_33_22;
    wire token_33_22;
    wire dep_chan_vld_34_22;
    wire [34:0] dep_chan_data_34_22;
    wire token_34_22;
    wire [16:0] proc_23_data_FIFO_blk;
    wire [16:0] proc_23_data_PIPO_blk;
    wire [16:0] proc_23_start_FIFO_blk;
    wire [16:0] proc_23_TLF_FIFO_blk;
    wire [16:0] proc_23_input_sync_blk;
    wire [16:0] proc_23_output_sync_blk;
    wire [16:0] proc_dep_vld_vec_23;
    reg [16:0] proc_dep_vld_vec_23_reg;
    wire [16:0] in_chan_dep_vld_vec_23;
    wire [594:0] in_chan_dep_data_vec_23;
    wire [16:0] token_in_vec_23;
    wire [16:0] out_chan_dep_vld_vec_23;
    wire [34:0] out_chan_dep_data_23;
    wire [16:0] token_out_vec_23;
    wire dl_detect_out_23;
    wire dep_chan_vld_0_23;
    wire [34:0] dep_chan_data_0_23;
    wire token_0_23;
    wire dep_chan_vld_7_23;
    wire [34:0] dep_chan_data_7_23;
    wire token_7_23;
    wire dep_chan_vld_19_23;
    wire [34:0] dep_chan_data_19_23;
    wire token_19_23;
    wire dep_chan_vld_20_23;
    wire [34:0] dep_chan_data_20_23;
    wire token_20_23;
    wire dep_chan_vld_21_23;
    wire [34:0] dep_chan_data_21_23;
    wire token_21_23;
    wire dep_chan_vld_22_23;
    wire [34:0] dep_chan_data_22_23;
    wire token_22_23;
    wire dep_chan_vld_24_23;
    wire [34:0] dep_chan_data_24_23;
    wire token_24_23;
    wire dep_chan_vld_25_23;
    wire [34:0] dep_chan_data_25_23;
    wire token_25_23;
    wire dep_chan_vld_26_23;
    wire [34:0] dep_chan_data_26_23;
    wire token_26_23;
    wire dep_chan_vld_27_23;
    wire [34:0] dep_chan_data_27_23;
    wire token_27_23;
    wire dep_chan_vld_28_23;
    wire [34:0] dep_chan_data_28_23;
    wire token_28_23;
    wire dep_chan_vld_29_23;
    wire [34:0] dep_chan_data_29_23;
    wire token_29_23;
    wire dep_chan_vld_30_23;
    wire [34:0] dep_chan_data_30_23;
    wire token_30_23;
    wire dep_chan_vld_31_23;
    wire [34:0] dep_chan_data_31_23;
    wire token_31_23;
    wire dep_chan_vld_32_23;
    wire [34:0] dep_chan_data_32_23;
    wire token_32_23;
    wire dep_chan_vld_33_23;
    wire [34:0] dep_chan_data_33_23;
    wire token_33_23;
    wire dep_chan_vld_34_23;
    wire [34:0] dep_chan_data_34_23;
    wire token_34_23;
    wire [16:0] proc_24_data_FIFO_blk;
    wire [16:0] proc_24_data_PIPO_blk;
    wire [16:0] proc_24_start_FIFO_blk;
    wire [16:0] proc_24_TLF_FIFO_blk;
    wire [16:0] proc_24_input_sync_blk;
    wire [16:0] proc_24_output_sync_blk;
    wire [16:0] proc_dep_vld_vec_24;
    reg [16:0] proc_dep_vld_vec_24_reg;
    wire [16:0] in_chan_dep_vld_vec_24;
    wire [594:0] in_chan_dep_data_vec_24;
    wire [16:0] token_in_vec_24;
    wire [16:0] out_chan_dep_vld_vec_24;
    wire [34:0] out_chan_dep_data_24;
    wire [16:0] token_out_vec_24;
    wire dl_detect_out_24;
    wire dep_chan_vld_0_24;
    wire [34:0] dep_chan_data_0_24;
    wire token_0_24;
    wire dep_chan_vld_8_24;
    wire [34:0] dep_chan_data_8_24;
    wire token_8_24;
    wire dep_chan_vld_19_24;
    wire [34:0] dep_chan_data_19_24;
    wire token_19_24;
    wire dep_chan_vld_20_24;
    wire [34:0] dep_chan_data_20_24;
    wire token_20_24;
    wire dep_chan_vld_21_24;
    wire [34:0] dep_chan_data_21_24;
    wire token_21_24;
    wire dep_chan_vld_22_24;
    wire [34:0] dep_chan_data_22_24;
    wire token_22_24;
    wire dep_chan_vld_23_24;
    wire [34:0] dep_chan_data_23_24;
    wire token_23_24;
    wire dep_chan_vld_25_24;
    wire [34:0] dep_chan_data_25_24;
    wire token_25_24;
    wire dep_chan_vld_26_24;
    wire [34:0] dep_chan_data_26_24;
    wire token_26_24;
    wire dep_chan_vld_27_24;
    wire [34:0] dep_chan_data_27_24;
    wire token_27_24;
    wire dep_chan_vld_28_24;
    wire [34:0] dep_chan_data_28_24;
    wire token_28_24;
    wire dep_chan_vld_29_24;
    wire [34:0] dep_chan_data_29_24;
    wire token_29_24;
    wire dep_chan_vld_30_24;
    wire [34:0] dep_chan_data_30_24;
    wire token_30_24;
    wire dep_chan_vld_31_24;
    wire [34:0] dep_chan_data_31_24;
    wire token_31_24;
    wire dep_chan_vld_32_24;
    wire [34:0] dep_chan_data_32_24;
    wire token_32_24;
    wire dep_chan_vld_33_24;
    wire [34:0] dep_chan_data_33_24;
    wire token_33_24;
    wire dep_chan_vld_34_24;
    wire [34:0] dep_chan_data_34_24;
    wire token_34_24;
    wire [16:0] proc_25_data_FIFO_blk;
    wire [16:0] proc_25_data_PIPO_blk;
    wire [16:0] proc_25_start_FIFO_blk;
    wire [16:0] proc_25_TLF_FIFO_blk;
    wire [16:0] proc_25_input_sync_blk;
    wire [16:0] proc_25_output_sync_blk;
    wire [16:0] proc_dep_vld_vec_25;
    reg [16:0] proc_dep_vld_vec_25_reg;
    wire [16:0] in_chan_dep_vld_vec_25;
    wire [594:0] in_chan_dep_data_vec_25;
    wire [16:0] token_in_vec_25;
    wire [16:0] out_chan_dep_vld_vec_25;
    wire [34:0] out_chan_dep_data_25;
    wire [16:0] token_out_vec_25;
    wire dl_detect_out_25;
    wire dep_chan_vld_0_25;
    wire [34:0] dep_chan_data_0_25;
    wire token_0_25;
    wire dep_chan_vld_9_25;
    wire [34:0] dep_chan_data_9_25;
    wire token_9_25;
    wire dep_chan_vld_19_25;
    wire [34:0] dep_chan_data_19_25;
    wire token_19_25;
    wire dep_chan_vld_20_25;
    wire [34:0] dep_chan_data_20_25;
    wire token_20_25;
    wire dep_chan_vld_21_25;
    wire [34:0] dep_chan_data_21_25;
    wire token_21_25;
    wire dep_chan_vld_22_25;
    wire [34:0] dep_chan_data_22_25;
    wire token_22_25;
    wire dep_chan_vld_23_25;
    wire [34:0] dep_chan_data_23_25;
    wire token_23_25;
    wire dep_chan_vld_24_25;
    wire [34:0] dep_chan_data_24_25;
    wire token_24_25;
    wire dep_chan_vld_26_25;
    wire [34:0] dep_chan_data_26_25;
    wire token_26_25;
    wire dep_chan_vld_27_25;
    wire [34:0] dep_chan_data_27_25;
    wire token_27_25;
    wire dep_chan_vld_28_25;
    wire [34:0] dep_chan_data_28_25;
    wire token_28_25;
    wire dep_chan_vld_29_25;
    wire [34:0] dep_chan_data_29_25;
    wire token_29_25;
    wire dep_chan_vld_30_25;
    wire [34:0] dep_chan_data_30_25;
    wire token_30_25;
    wire dep_chan_vld_31_25;
    wire [34:0] dep_chan_data_31_25;
    wire token_31_25;
    wire dep_chan_vld_32_25;
    wire [34:0] dep_chan_data_32_25;
    wire token_32_25;
    wire dep_chan_vld_33_25;
    wire [34:0] dep_chan_data_33_25;
    wire token_33_25;
    wire dep_chan_vld_34_25;
    wire [34:0] dep_chan_data_34_25;
    wire token_34_25;
    wire [16:0] proc_26_data_FIFO_blk;
    wire [16:0] proc_26_data_PIPO_blk;
    wire [16:0] proc_26_start_FIFO_blk;
    wire [16:0] proc_26_TLF_FIFO_blk;
    wire [16:0] proc_26_input_sync_blk;
    wire [16:0] proc_26_output_sync_blk;
    wire [16:0] proc_dep_vld_vec_26;
    reg [16:0] proc_dep_vld_vec_26_reg;
    wire [16:0] in_chan_dep_vld_vec_26;
    wire [594:0] in_chan_dep_data_vec_26;
    wire [16:0] token_in_vec_26;
    wire [16:0] out_chan_dep_vld_vec_26;
    wire [34:0] out_chan_dep_data_26;
    wire [16:0] token_out_vec_26;
    wire dl_detect_out_26;
    wire dep_chan_vld_0_26;
    wire [34:0] dep_chan_data_0_26;
    wire token_0_26;
    wire dep_chan_vld_10_26;
    wire [34:0] dep_chan_data_10_26;
    wire token_10_26;
    wire dep_chan_vld_19_26;
    wire [34:0] dep_chan_data_19_26;
    wire token_19_26;
    wire dep_chan_vld_20_26;
    wire [34:0] dep_chan_data_20_26;
    wire token_20_26;
    wire dep_chan_vld_21_26;
    wire [34:0] dep_chan_data_21_26;
    wire token_21_26;
    wire dep_chan_vld_22_26;
    wire [34:0] dep_chan_data_22_26;
    wire token_22_26;
    wire dep_chan_vld_23_26;
    wire [34:0] dep_chan_data_23_26;
    wire token_23_26;
    wire dep_chan_vld_24_26;
    wire [34:0] dep_chan_data_24_26;
    wire token_24_26;
    wire dep_chan_vld_25_26;
    wire [34:0] dep_chan_data_25_26;
    wire token_25_26;
    wire dep_chan_vld_27_26;
    wire [34:0] dep_chan_data_27_26;
    wire token_27_26;
    wire dep_chan_vld_28_26;
    wire [34:0] dep_chan_data_28_26;
    wire token_28_26;
    wire dep_chan_vld_29_26;
    wire [34:0] dep_chan_data_29_26;
    wire token_29_26;
    wire dep_chan_vld_30_26;
    wire [34:0] dep_chan_data_30_26;
    wire token_30_26;
    wire dep_chan_vld_31_26;
    wire [34:0] dep_chan_data_31_26;
    wire token_31_26;
    wire dep_chan_vld_32_26;
    wire [34:0] dep_chan_data_32_26;
    wire token_32_26;
    wire dep_chan_vld_33_26;
    wire [34:0] dep_chan_data_33_26;
    wire token_33_26;
    wire dep_chan_vld_34_26;
    wire [34:0] dep_chan_data_34_26;
    wire token_34_26;
    wire [16:0] proc_27_data_FIFO_blk;
    wire [16:0] proc_27_data_PIPO_blk;
    wire [16:0] proc_27_start_FIFO_blk;
    wire [16:0] proc_27_TLF_FIFO_blk;
    wire [16:0] proc_27_input_sync_blk;
    wire [16:0] proc_27_output_sync_blk;
    wire [16:0] proc_dep_vld_vec_27;
    reg [16:0] proc_dep_vld_vec_27_reg;
    wire [16:0] in_chan_dep_vld_vec_27;
    wire [594:0] in_chan_dep_data_vec_27;
    wire [16:0] token_in_vec_27;
    wire [16:0] out_chan_dep_vld_vec_27;
    wire [34:0] out_chan_dep_data_27;
    wire [16:0] token_out_vec_27;
    wire dl_detect_out_27;
    wire dep_chan_vld_0_27;
    wire [34:0] dep_chan_data_0_27;
    wire token_0_27;
    wire dep_chan_vld_11_27;
    wire [34:0] dep_chan_data_11_27;
    wire token_11_27;
    wire dep_chan_vld_19_27;
    wire [34:0] dep_chan_data_19_27;
    wire token_19_27;
    wire dep_chan_vld_20_27;
    wire [34:0] dep_chan_data_20_27;
    wire token_20_27;
    wire dep_chan_vld_21_27;
    wire [34:0] dep_chan_data_21_27;
    wire token_21_27;
    wire dep_chan_vld_22_27;
    wire [34:0] dep_chan_data_22_27;
    wire token_22_27;
    wire dep_chan_vld_23_27;
    wire [34:0] dep_chan_data_23_27;
    wire token_23_27;
    wire dep_chan_vld_24_27;
    wire [34:0] dep_chan_data_24_27;
    wire token_24_27;
    wire dep_chan_vld_25_27;
    wire [34:0] dep_chan_data_25_27;
    wire token_25_27;
    wire dep_chan_vld_26_27;
    wire [34:0] dep_chan_data_26_27;
    wire token_26_27;
    wire dep_chan_vld_28_27;
    wire [34:0] dep_chan_data_28_27;
    wire token_28_27;
    wire dep_chan_vld_29_27;
    wire [34:0] dep_chan_data_29_27;
    wire token_29_27;
    wire dep_chan_vld_30_27;
    wire [34:0] dep_chan_data_30_27;
    wire token_30_27;
    wire dep_chan_vld_31_27;
    wire [34:0] dep_chan_data_31_27;
    wire token_31_27;
    wire dep_chan_vld_32_27;
    wire [34:0] dep_chan_data_32_27;
    wire token_32_27;
    wire dep_chan_vld_33_27;
    wire [34:0] dep_chan_data_33_27;
    wire token_33_27;
    wire dep_chan_vld_34_27;
    wire [34:0] dep_chan_data_34_27;
    wire token_34_27;
    wire [16:0] proc_28_data_FIFO_blk;
    wire [16:0] proc_28_data_PIPO_blk;
    wire [16:0] proc_28_start_FIFO_blk;
    wire [16:0] proc_28_TLF_FIFO_blk;
    wire [16:0] proc_28_input_sync_blk;
    wire [16:0] proc_28_output_sync_blk;
    wire [16:0] proc_dep_vld_vec_28;
    reg [16:0] proc_dep_vld_vec_28_reg;
    wire [16:0] in_chan_dep_vld_vec_28;
    wire [594:0] in_chan_dep_data_vec_28;
    wire [16:0] token_in_vec_28;
    wire [16:0] out_chan_dep_vld_vec_28;
    wire [34:0] out_chan_dep_data_28;
    wire [16:0] token_out_vec_28;
    wire dl_detect_out_28;
    wire dep_chan_vld_0_28;
    wire [34:0] dep_chan_data_0_28;
    wire token_0_28;
    wire dep_chan_vld_12_28;
    wire [34:0] dep_chan_data_12_28;
    wire token_12_28;
    wire dep_chan_vld_19_28;
    wire [34:0] dep_chan_data_19_28;
    wire token_19_28;
    wire dep_chan_vld_20_28;
    wire [34:0] dep_chan_data_20_28;
    wire token_20_28;
    wire dep_chan_vld_21_28;
    wire [34:0] dep_chan_data_21_28;
    wire token_21_28;
    wire dep_chan_vld_22_28;
    wire [34:0] dep_chan_data_22_28;
    wire token_22_28;
    wire dep_chan_vld_23_28;
    wire [34:0] dep_chan_data_23_28;
    wire token_23_28;
    wire dep_chan_vld_24_28;
    wire [34:0] dep_chan_data_24_28;
    wire token_24_28;
    wire dep_chan_vld_25_28;
    wire [34:0] dep_chan_data_25_28;
    wire token_25_28;
    wire dep_chan_vld_26_28;
    wire [34:0] dep_chan_data_26_28;
    wire token_26_28;
    wire dep_chan_vld_27_28;
    wire [34:0] dep_chan_data_27_28;
    wire token_27_28;
    wire dep_chan_vld_29_28;
    wire [34:0] dep_chan_data_29_28;
    wire token_29_28;
    wire dep_chan_vld_30_28;
    wire [34:0] dep_chan_data_30_28;
    wire token_30_28;
    wire dep_chan_vld_31_28;
    wire [34:0] dep_chan_data_31_28;
    wire token_31_28;
    wire dep_chan_vld_32_28;
    wire [34:0] dep_chan_data_32_28;
    wire token_32_28;
    wire dep_chan_vld_33_28;
    wire [34:0] dep_chan_data_33_28;
    wire token_33_28;
    wire dep_chan_vld_34_28;
    wire [34:0] dep_chan_data_34_28;
    wire token_34_28;
    wire [16:0] proc_29_data_FIFO_blk;
    wire [16:0] proc_29_data_PIPO_blk;
    wire [16:0] proc_29_start_FIFO_blk;
    wire [16:0] proc_29_TLF_FIFO_blk;
    wire [16:0] proc_29_input_sync_blk;
    wire [16:0] proc_29_output_sync_blk;
    wire [16:0] proc_dep_vld_vec_29;
    reg [16:0] proc_dep_vld_vec_29_reg;
    wire [16:0] in_chan_dep_vld_vec_29;
    wire [594:0] in_chan_dep_data_vec_29;
    wire [16:0] token_in_vec_29;
    wire [16:0] out_chan_dep_vld_vec_29;
    wire [34:0] out_chan_dep_data_29;
    wire [16:0] token_out_vec_29;
    wire dl_detect_out_29;
    wire dep_chan_vld_0_29;
    wire [34:0] dep_chan_data_0_29;
    wire token_0_29;
    wire dep_chan_vld_13_29;
    wire [34:0] dep_chan_data_13_29;
    wire token_13_29;
    wire dep_chan_vld_19_29;
    wire [34:0] dep_chan_data_19_29;
    wire token_19_29;
    wire dep_chan_vld_20_29;
    wire [34:0] dep_chan_data_20_29;
    wire token_20_29;
    wire dep_chan_vld_21_29;
    wire [34:0] dep_chan_data_21_29;
    wire token_21_29;
    wire dep_chan_vld_22_29;
    wire [34:0] dep_chan_data_22_29;
    wire token_22_29;
    wire dep_chan_vld_23_29;
    wire [34:0] dep_chan_data_23_29;
    wire token_23_29;
    wire dep_chan_vld_24_29;
    wire [34:0] dep_chan_data_24_29;
    wire token_24_29;
    wire dep_chan_vld_25_29;
    wire [34:0] dep_chan_data_25_29;
    wire token_25_29;
    wire dep_chan_vld_26_29;
    wire [34:0] dep_chan_data_26_29;
    wire token_26_29;
    wire dep_chan_vld_27_29;
    wire [34:0] dep_chan_data_27_29;
    wire token_27_29;
    wire dep_chan_vld_28_29;
    wire [34:0] dep_chan_data_28_29;
    wire token_28_29;
    wire dep_chan_vld_30_29;
    wire [34:0] dep_chan_data_30_29;
    wire token_30_29;
    wire dep_chan_vld_31_29;
    wire [34:0] dep_chan_data_31_29;
    wire token_31_29;
    wire dep_chan_vld_32_29;
    wire [34:0] dep_chan_data_32_29;
    wire token_32_29;
    wire dep_chan_vld_33_29;
    wire [34:0] dep_chan_data_33_29;
    wire token_33_29;
    wire dep_chan_vld_34_29;
    wire [34:0] dep_chan_data_34_29;
    wire token_34_29;
    wire [16:0] proc_30_data_FIFO_blk;
    wire [16:0] proc_30_data_PIPO_blk;
    wire [16:0] proc_30_start_FIFO_blk;
    wire [16:0] proc_30_TLF_FIFO_blk;
    wire [16:0] proc_30_input_sync_blk;
    wire [16:0] proc_30_output_sync_blk;
    wire [16:0] proc_dep_vld_vec_30;
    reg [16:0] proc_dep_vld_vec_30_reg;
    wire [16:0] in_chan_dep_vld_vec_30;
    wire [594:0] in_chan_dep_data_vec_30;
    wire [16:0] token_in_vec_30;
    wire [16:0] out_chan_dep_vld_vec_30;
    wire [34:0] out_chan_dep_data_30;
    wire [16:0] token_out_vec_30;
    wire dl_detect_out_30;
    wire dep_chan_vld_0_30;
    wire [34:0] dep_chan_data_0_30;
    wire token_0_30;
    wire dep_chan_vld_14_30;
    wire [34:0] dep_chan_data_14_30;
    wire token_14_30;
    wire dep_chan_vld_19_30;
    wire [34:0] dep_chan_data_19_30;
    wire token_19_30;
    wire dep_chan_vld_20_30;
    wire [34:0] dep_chan_data_20_30;
    wire token_20_30;
    wire dep_chan_vld_21_30;
    wire [34:0] dep_chan_data_21_30;
    wire token_21_30;
    wire dep_chan_vld_22_30;
    wire [34:0] dep_chan_data_22_30;
    wire token_22_30;
    wire dep_chan_vld_23_30;
    wire [34:0] dep_chan_data_23_30;
    wire token_23_30;
    wire dep_chan_vld_24_30;
    wire [34:0] dep_chan_data_24_30;
    wire token_24_30;
    wire dep_chan_vld_25_30;
    wire [34:0] dep_chan_data_25_30;
    wire token_25_30;
    wire dep_chan_vld_26_30;
    wire [34:0] dep_chan_data_26_30;
    wire token_26_30;
    wire dep_chan_vld_27_30;
    wire [34:0] dep_chan_data_27_30;
    wire token_27_30;
    wire dep_chan_vld_28_30;
    wire [34:0] dep_chan_data_28_30;
    wire token_28_30;
    wire dep_chan_vld_29_30;
    wire [34:0] dep_chan_data_29_30;
    wire token_29_30;
    wire dep_chan_vld_31_30;
    wire [34:0] dep_chan_data_31_30;
    wire token_31_30;
    wire dep_chan_vld_32_30;
    wire [34:0] dep_chan_data_32_30;
    wire token_32_30;
    wire dep_chan_vld_33_30;
    wire [34:0] dep_chan_data_33_30;
    wire token_33_30;
    wire dep_chan_vld_34_30;
    wire [34:0] dep_chan_data_34_30;
    wire token_34_30;
    wire [16:0] proc_31_data_FIFO_blk;
    wire [16:0] proc_31_data_PIPO_blk;
    wire [16:0] proc_31_start_FIFO_blk;
    wire [16:0] proc_31_TLF_FIFO_blk;
    wire [16:0] proc_31_input_sync_blk;
    wire [16:0] proc_31_output_sync_blk;
    wire [16:0] proc_dep_vld_vec_31;
    reg [16:0] proc_dep_vld_vec_31_reg;
    wire [16:0] in_chan_dep_vld_vec_31;
    wire [594:0] in_chan_dep_data_vec_31;
    wire [16:0] token_in_vec_31;
    wire [16:0] out_chan_dep_vld_vec_31;
    wire [34:0] out_chan_dep_data_31;
    wire [16:0] token_out_vec_31;
    wire dl_detect_out_31;
    wire dep_chan_vld_0_31;
    wire [34:0] dep_chan_data_0_31;
    wire token_0_31;
    wire dep_chan_vld_15_31;
    wire [34:0] dep_chan_data_15_31;
    wire token_15_31;
    wire dep_chan_vld_19_31;
    wire [34:0] dep_chan_data_19_31;
    wire token_19_31;
    wire dep_chan_vld_20_31;
    wire [34:0] dep_chan_data_20_31;
    wire token_20_31;
    wire dep_chan_vld_21_31;
    wire [34:0] dep_chan_data_21_31;
    wire token_21_31;
    wire dep_chan_vld_22_31;
    wire [34:0] dep_chan_data_22_31;
    wire token_22_31;
    wire dep_chan_vld_23_31;
    wire [34:0] dep_chan_data_23_31;
    wire token_23_31;
    wire dep_chan_vld_24_31;
    wire [34:0] dep_chan_data_24_31;
    wire token_24_31;
    wire dep_chan_vld_25_31;
    wire [34:0] dep_chan_data_25_31;
    wire token_25_31;
    wire dep_chan_vld_26_31;
    wire [34:0] dep_chan_data_26_31;
    wire token_26_31;
    wire dep_chan_vld_27_31;
    wire [34:0] dep_chan_data_27_31;
    wire token_27_31;
    wire dep_chan_vld_28_31;
    wire [34:0] dep_chan_data_28_31;
    wire token_28_31;
    wire dep_chan_vld_29_31;
    wire [34:0] dep_chan_data_29_31;
    wire token_29_31;
    wire dep_chan_vld_30_31;
    wire [34:0] dep_chan_data_30_31;
    wire token_30_31;
    wire dep_chan_vld_32_31;
    wire [34:0] dep_chan_data_32_31;
    wire token_32_31;
    wire dep_chan_vld_33_31;
    wire [34:0] dep_chan_data_33_31;
    wire token_33_31;
    wire dep_chan_vld_34_31;
    wire [34:0] dep_chan_data_34_31;
    wire token_34_31;
    wire [16:0] proc_32_data_FIFO_blk;
    wire [16:0] proc_32_data_PIPO_blk;
    wire [16:0] proc_32_start_FIFO_blk;
    wire [16:0] proc_32_TLF_FIFO_blk;
    wire [16:0] proc_32_input_sync_blk;
    wire [16:0] proc_32_output_sync_blk;
    wire [16:0] proc_dep_vld_vec_32;
    reg [16:0] proc_dep_vld_vec_32_reg;
    wire [16:0] in_chan_dep_vld_vec_32;
    wire [594:0] in_chan_dep_data_vec_32;
    wire [16:0] token_in_vec_32;
    wire [16:0] out_chan_dep_vld_vec_32;
    wire [34:0] out_chan_dep_data_32;
    wire [16:0] token_out_vec_32;
    wire dl_detect_out_32;
    wire dep_chan_vld_0_32;
    wire [34:0] dep_chan_data_0_32;
    wire token_0_32;
    wire dep_chan_vld_16_32;
    wire [34:0] dep_chan_data_16_32;
    wire token_16_32;
    wire dep_chan_vld_19_32;
    wire [34:0] dep_chan_data_19_32;
    wire token_19_32;
    wire dep_chan_vld_20_32;
    wire [34:0] dep_chan_data_20_32;
    wire token_20_32;
    wire dep_chan_vld_21_32;
    wire [34:0] dep_chan_data_21_32;
    wire token_21_32;
    wire dep_chan_vld_22_32;
    wire [34:0] dep_chan_data_22_32;
    wire token_22_32;
    wire dep_chan_vld_23_32;
    wire [34:0] dep_chan_data_23_32;
    wire token_23_32;
    wire dep_chan_vld_24_32;
    wire [34:0] dep_chan_data_24_32;
    wire token_24_32;
    wire dep_chan_vld_25_32;
    wire [34:0] dep_chan_data_25_32;
    wire token_25_32;
    wire dep_chan_vld_26_32;
    wire [34:0] dep_chan_data_26_32;
    wire token_26_32;
    wire dep_chan_vld_27_32;
    wire [34:0] dep_chan_data_27_32;
    wire token_27_32;
    wire dep_chan_vld_28_32;
    wire [34:0] dep_chan_data_28_32;
    wire token_28_32;
    wire dep_chan_vld_29_32;
    wire [34:0] dep_chan_data_29_32;
    wire token_29_32;
    wire dep_chan_vld_30_32;
    wire [34:0] dep_chan_data_30_32;
    wire token_30_32;
    wire dep_chan_vld_31_32;
    wire [34:0] dep_chan_data_31_32;
    wire token_31_32;
    wire dep_chan_vld_33_32;
    wire [34:0] dep_chan_data_33_32;
    wire token_33_32;
    wire dep_chan_vld_34_32;
    wire [34:0] dep_chan_data_34_32;
    wire token_34_32;
    wire [16:0] proc_33_data_FIFO_blk;
    wire [16:0] proc_33_data_PIPO_blk;
    wire [16:0] proc_33_start_FIFO_blk;
    wire [16:0] proc_33_TLF_FIFO_blk;
    wire [16:0] proc_33_input_sync_blk;
    wire [16:0] proc_33_output_sync_blk;
    wire [16:0] proc_dep_vld_vec_33;
    reg [16:0] proc_dep_vld_vec_33_reg;
    wire [16:0] in_chan_dep_vld_vec_33;
    wire [594:0] in_chan_dep_data_vec_33;
    wire [16:0] token_in_vec_33;
    wire [16:0] out_chan_dep_vld_vec_33;
    wire [34:0] out_chan_dep_data_33;
    wire [16:0] token_out_vec_33;
    wire dl_detect_out_33;
    wire dep_chan_vld_0_33;
    wire [34:0] dep_chan_data_0_33;
    wire token_0_33;
    wire dep_chan_vld_17_33;
    wire [34:0] dep_chan_data_17_33;
    wire token_17_33;
    wire dep_chan_vld_19_33;
    wire [34:0] dep_chan_data_19_33;
    wire token_19_33;
    wire dep_chan_vld_20_33;
    wire [34:0] dep_chan_data_20_33;
    wire token_20_33;
    wire dep_chan_vld_21_33;
    wire [34:0] dep_chan_data_21_33;
    wire token_21_33;
    wire dep_chan_vld_22_33;
    wire [34:0] dep_chan_data_22_33;
    wire token_22_33;
    wire dep_chan_vld_23_33;
    wire [34:0] dep_chan_data_23_33;
    wire token_23_33;
    wire dep_chan_vld_24_33;
    wire [34:0] dep_chan_data_24_33;
    wire token_24_33;
    wire dep_chan_vld_25_33;
    wire [34:0] dep_chan_data_25_33;
    wire token_25_33;
    wire dep_chan_vld_26_33;
    wire [34:0] dep_chan_data_26_33;
    wire token_26_33;
    wire dep_chan_vld_27_33;
    wire [34:0] dep_chan_data_27_33;
    wire token_27_33;
    wire dep_chan_vld_28_33;
    wire [34:0] dep_chan_data_28_33;
    wire token_28_33;
    wire dep_chan_vld_29_33;
    wire [34:0] dep_chan_data_29_33;
    wire token_29_33;
    wire dep_chan_vld_30_33;
    wire [34:0] dep_chan_data_30_33;
    wire token_30_33;
    wire dep_chan_vld_31_33;
    wire [34:0] dep_chan_data_31_33;
    wire token_31_33;
    wire dep_chan_vld_32_33;
    wire [34:0] dep_chan_data_32_33;
    wire token_32_33;
    wire dep_chan_vld_34_33;
    wire [34:0] dep_chan_data_34_33;
    wire token_34_33;
    wire [16:0] proc_34_data_FIFO_blk;
    wire [16:0] proc_34_data_PIPO_blk;
    wire [16:0] proc_34_start_FIFO_blk;
    wire [16:0] proc_34_TLF_FIFO_blk;
    wire [16:0] proc_34_input_sync_blk;
    wire [16:0] proc_34_output_sync_blk;
    wire [16:0] proc_dep_vld_vec_34;
    reg [16:0] proc_dep_vld_vec_34_reg;
    wire [16:0] in_chan_dep_vld_vec_34;
    wire [594:0] in_chan_dep_data_vec_34;
    wire [16:0] token_in_vec_34;
    wire [16:0] out_chan_dep_vld_vec_34;
    wire [34:0] out_chan_dep_data_34;
    wire [16:0] token_out_vec_34;
    wire dl_detect_out_34;
    wire dep_chan_vld_0_34;
    wire [34:0] dep_chan_data_0_34;
    wire token_0_34;
    wire dep_chan_vld_18_34;
    wire [34:0] dep_chan_data_18_34;
    wire token_18_34;
    wire dep_chan_vld_19_34;
    wire [34:0] dep_chan_data_19_34;
    wire token_19_34;
    wire dep_chan_vld_20_34;
    wire [34:0] dep_chan_data_20_34;
    wire token_20_34;
    wire dep_chan_vld_21_34;
    wire [34:0] dep_chan_data_21_34;
    wire token_21_34;
    wire dep_chan_vld_22_34;
    wire [34:0] dep_chan_data_22_34;
    wire token_22_34;
    wire dep_chan_vld_23_34;
    wire [34:0] dep_chan_data_23_34;
    wire token_23_34;
    wire dep_chan_vld_24_34;
    wire [34:0] dep_chan_data_24_34;
    wire token_24_34;
    wire dep_chan_vld_25_34;
    wire [34:0] dep_chan_data_25_34;
    wire token_25_34;
    wire dep_chan_vld_26_34;
    wire [34:0] dep_chan_data_26_34;
    wire token_26_34;
    wire dep_chan_vld_27_34;
    wire [34:0] dep_chan_data_27_34;
    wire token_27_34;
    wire dep_chan_vld_28_34;
    wire [34:0] dep_chan_data_28_34;
    wire token_28_34;
    wire dep_chan_vld_29_34;
    wire [34:0] dep_chan_data_29_34;
    wire token_29_34;
    wire dep_chan_vld_30_34;
    wire [34:0] dep_chan_data_30_34;
    wire token_30_34;
    wire dep_chan_vld_31_34;
    wire [34:0] dep_chan_data_31_34;
    wire token_31_34;
    wire dep_chan_vld_32_34;
    wire [34:0] dep_chan_data_32_34;
    wire token_32_34;
    wire dep_chan_vld_33_34;
    wire [34:0] dep_chan_data_33_34;
    wire token_33_34;
    wire [34:0] dl_in_vec;
    wire dl_detect_out;
    wire token_clear;
    reg [34:0] origin;

    reg ap_done_reg_0;// for module write_back48_U0
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_0 <= 'b0;
        end
        else begin
            ap_done_reg_0 <= write_back48_U0.ap_done & ~write_back48_U0.ap_continue;
        end
    end

    reg ap_done_reg_1;// for module write_back49_U0
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_1 <= 'b0;
        end
        else begin
            ap_done_reg_1 <= write_back49_U0.ap_done & ~write_back49_U0.ap_continue;
        end
    end

    reg ap_done_reg_2;// for module write_back50_U0
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_2 <= 'b0;
        end
        else begin
            ap_done_reg_2 <= write_back50_U0.ap_done & ~write_back50_U0.ap_continue;
        end
    end

    reg ap_done_reg_3;// for module write_back51_U0
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_3 <= 'b0;
        end
        else begin
            ap_done_reg_3 <= write_back51_U0.ap_done & ~write_back51_U0.ap_continue;
        end
    end

    reg ap_done_reg_4;// for module write_back52_U0
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_4 <= 'b0;
        end
        else begin
            ap_done_reg_4 <= write_back52_U0.ap_done & ~write_back52_U0.ap_continue;
        end
    end

    reg ap_done_reg_5;// for module write_back53_U0
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_5 <= 'b0;
        end
        else begin
            ap_done_reg_5 <= write_back53_U0.ap_done & ~write_back53_U0.ap_continue;
        end
    end

    reg ap_done_reg_6;// for module write_back54_U0
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_6 <= 'b0;
        end
        else begin
            ap_done_reg_6 <= write_back54_U0.ap_done & ~write_back54_U0.ap_continue;
        end
    end

    reg ap_done_reg_7;// for module write_back55_U0
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_7 <= 'b0;
        end
        else begin
            ap_done_reg_7 <= write_back55_U0.ap_done & ~write_back55_U0.ap_continue;
        end
    end

    reg ap_done_reg_8;// for module write_back56_U0
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_8 <= 'b0;
        end
        else begin
            ap_done_reg_8 <= write_back56_U0.ap_done & ~write_back56_U0.ap_continue;
        end
    end

    reg ap_done_reg_9;// for module write_back57_U0
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_9 <= 'b0;
        end
        else begin
            ap_done_reg_9 <= write_back57_U0.ap_done & ~write_back57_U0.ap_continue;
        end
    end

    reg ap_done_reg_10;// for module write_back58_U0
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_10 <= 'b0;
        end
        else begin
            ap_done_reg_10 <= write_back58_U0.ap_done & ~write_back58_U0.ap_continue;
        end
    end

    reg ap_done_reg_11;// for module write_back59_U0
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_11 <= 'b0;
        end
        else begin
            ap_done_reg_11 <= write_back59_U0.ap_done & ~write_back59_U0.ap_continue;
        end
    end

    reg ap_done_reg_12;// for module write_back60_U0
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_12 <= 'b0;
        end
        else begin
            ap_done_reg_12 <= write_back60_U0.ap_done & ~write_back60_U0.ap_continue;
        end
    end

    reg ap_done_reg_13;// for module write_back61_U0
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_13 <= 'b0;
        end
        else begin
            ap_done_reg_13 <= write_back61_U0.ap_done & ~write_back61_U0.ap_continue;
        end
    end

    reg ap_done_reg_14;// for module write_back62_U0
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_14 <= 'b0;
        end
        else begin
            ap_done_reg_14 <= write_back62_U0.ap_done & ~write_back62_U0.ap_continue;
        end
    end

    reg ap_done_reg_15;// for module write_back63_U0
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            ap_done_reg_15 <= 'b0;
        end
        else begin
            ap_done_reg_15 <= write_back63_U0.ap_done & ~write_back63_U0.ap_continue;
        end
    end

reg [15:0] trans_in_cnt_0;// for process kernel_pr_entry98_U0
always @(negedge reset or posedge clock) begin
    if (~reset) begin
         trans_in_cnt_0 <= 16'h0;
    end
    else if (kernel_pr_entry98_U0.start_write == 1'b1) begin
        trans_in_cnt_0 <= trans_in_cnt_0 + 16'h1;
    end
    else begin
        trans_in_cnt_0 <= trans_in_cnt_0;
    end
end

reg [15:0] trans_out_cnt_0;// for process kernel_pr_entry98_U0
always @(negedge reset or posedge clock) begin
    if (~reset) begin
         trans_out_cnt_0 <= 16'h0;
    end
    else if (kernel_pr_entry98_U0.ap_done == 1'b1 && kernel_pr_entry98_U0.ap_continue == 1'b1) begin
        trans_out_cnt_0 <= trans_out_cnt_0 + 16'h1;
    end
    else begin
        trans_out_cnt_0 <= trans_out_cnt_0;
    end
end

    // Process: kernel_pr_entry98_U0
    kernel_pr_hls_deadlock_detect_unit #(35, 0, 34, 34) kernel_pr_hls_deadlock_detect_unit_0 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_0),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_0),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_0),
        .token_in_vec(token_in_vec_0),
        .dl_detect_in(dl_detect_out),
        .origin(origin[0]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_0),
        .out_chan_dep_data(out_chan_dep_data_0),
        .token_out_vec(token_out_vec_0),
        .dl_detect_out(dl_in_vec[0]));

    assign proc_0_data_FIFO_blk[0] = 1'b0 | (~kernel_pr_entry98_U0.H_write0_out_blk_n) | (~kernel_pr_entry98_U0.hyperedge_size_out_blk_n);
    assign proc_0_data_PIPO_blk[0] = 1'b0;
    assign proc_0_start_FIFO_blk[0] = 1'b0 | (~start_for_write_back48_U0_U.if_full_n & kernel_pr_entry98_U0.ap_start & ~kernel_pr_entry98_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_write_back48_U0_U.if_read);
    assign proc_0_TLF_FIFO_blk[0] = 1'b0;
    assign proc_0_input_sync_blk[0] = 1'b0;
    assign proc_0_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_0[0] = dl_detect_out ? proc_dep_vld_vec_0_reg[0] : (proc_0_data_FIFO_blk[0] | proc_0_data_PIPO_blk[0] | proc_0_start_FIFO_blk[0] | proc_0_TLF_FIFO_blk[0] | proc_0_input_sync_blk[0] | proc_0_output_sync_blk[0]);
    assign proc_0_data_FIFO_blk[1] = 1'b0 | (~kernel_pr_entry98_U0.H_write1_out_blk_n) | (~kernel_pr_entry98_U0.hyperedge_size_out1_blk_n);
    assign proc_0_data_PIPO_blk[1] = 1'b0;
    assign proc_0_start_FIFO_blk[1] = 1'b0 | (~start_for_write_back49_U0_U.if_full_n & kernel_pr_entry98_U0.ap_start & ~kernel_pr_entry98_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_write_back49_U0_U.if_read);
    assign proc_0_TLF_FIFO_blk[1] = 1'b0;
    assign proc_0_input_sync_blk[1] = 1'b0;
    assign proc_0_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_0[1] = dl_detect_out ? proc_dep_vld_vec_0_reg[1] : (proc_0_data_FIFO_blk[1] | proc_0_data_PIPO_blk[1] | proc_0_start_FIFO_blk[1] | proc_0_TLF_FIFO_blk[1] | proc_0_input_sync_blk[1] | proc_0_output_sync_blk[1]);
    assign proc_0_data_FIFO_blk[2] = 1'b0 | (~kernel_pr_entry98_U0.H_write2_out_blk_n) | (~kernel_pr_entry98_U0.hyperedge_size_out2_blk_n);
    assign proc_0_data_PIPO_blk[2] = 1'b0;
    assign proc_0_start_FIFO_blk[2] = 1'b0 | (~start_for_write_back50_U0_U.if_full_n & kernel_pr_entry98_U0.ap_start & ~kernel_pr_entry98_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_write_back50_U0_U.if_read);
    assign proc_0_TLF_FIFO_blk[2] = 1'b0;
    assign proc_0_input_sync_blk[2] = 1'b0;
    assign proc_0_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_0[2] = dl_detect_out ? proc_dep_vld_vec_0_reg[2] : (proc_0_data_FIFO_blk[2] | proc_0_data_PIPO_blk[2] | proc_0_start_FIFO_blk[2] | proc_0_TLF_FIFO_blk[2] | proc_0_input_sync_blk[2] | proc_0_output_sync_blk[2]);
    assign proc_0_data_FIFO_blk[3] = 1'b0 | (~kernel_pr_entry98_U0.H_write3_out_blk_n) | (~kernel_pr_entry98_U0.hyperedge_size_out3_blk_n);
    assign proc_0_data_PIPO_blk[3] = 1'b0;
    assign proc_0_start_FIFO_blk[3] = 1'b0 | (~start_for_write_back51_U0_U.if_full_n & kernel_pr_entry98_U0.ap_start & ~kernel_pr_entry98_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_write_back51_U0_U.if_read);
    assign proc_0_TLF_FIFO_blk[3] = 1'b0;
    assign proc_0_input_sync_blk[3] = 1'b0;
    assign proc_0_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_0[3] = dl_detect_out ? proc_dep_vld_vec_0_reg[3] : (proc_0_data_FIFO_blk[3] | proc_0_data_PIPO_blk[3] | proc_0_start_FIFO_blk[3] | proc_0_TLF_FIFO_blk[3] | proc_0_input_sync_blk[3] | proc_0_output_sync_blk[3]);
    assign proc_0_data_FIFO_blk[4] = 1'b0 | (~kernel_pr_entry98_U0.H_write4_out_blk_n) | (~kernel_pr_entry98_U0.hyperedge_size_out4_blk_n);
    assign proc_0_data_PIPO_blk[4] = 1'b0;
    assign proc_0_start_FIFO_blk[4] = 1'b0 | (~start_for_write_back52_U0_U.if_full_n & kernel_pr_entry98_U0.ap_start & ~kernel_pr_entry98_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_write_back52_U0_U.if_read);
    assign proc_0_TLF_FIFO_blk[4] = 1'b0;
    assign proc_0_input_sync_blk[4] = 1'b0;
    assign proc_0_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_0[4] = dl_detect_out ? proc_dep_vld_vec_0_reg[4] : (proc_0_data_FIFO_blk[4] | proc_0_data_PIPO_blk[4] | proc_0_start_FIFO_blk[4] | proc_0_TLF_FIFO_blk[4] | proc_0_input_sync_blk[4] | proc_0_output_sync_blk[4]);
    assign proc_0_data_FIFO_blk[5] = 1'b0 | (~kernel_pr_entry98_U0.H_write5_out_blk_n) | (~kernel_pr_entry98_U0.hyperedge_size_out5_blk_n);
    assign proc_0_data_PIPO_blk[5] = 1'b0;
    assign proc_0_start_FIFO_blk[5] = 1'b0 | (~start_for_write_back53_U0_U.if_full_n & kernel_pr_entry98_U0.ap_start & ~kernel_pr_entry98_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_write_back53_U0_U.if_read);
    assign proc_0_TLF_FIFO_blk[5] = 1'b0;
    assign proc_0_input_sync_blk[5] = 1'b0;
    assign proc_0_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_0[5] = dl_detect_out ? proc_dep_vld_vec_0_reg[5] : (proc_0_data_FIFO_blk[5] | proc_0_data_PIPO_blk[5] | proc_0_start_FIFO_blk[5] | proc_0_TLF_FIFO_blk[5] | proc_0_input_sync_blk[5] | proc_0_output_sync_blk[5]);
    assign proc_0_data_FIFO_blk[6] = 1'b0 | (~kernel_pr_entry98_U0.H_write6_out_blk_n) | (~kernel_pr_entry98_U0.hyperedge_size_out6_blk_n);
    assign proc_0_data_PIPO_blk[6] = 1'b0;
    assign proc_0_start_FIFO_blk[6] = 1'b0 | (~start_for_write_back54_U0_U.if_full_n & kernel_pr_entry98_U0.ap_start & ~kernel_pr_entry98_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_write_back54_U0_U.if_read);
    assign proc_0_TLF_FIFO_blk[6] = 1'b0;
    assign proc_0_input_sync_blk[6] = 1'b0;
    assign proc_0_output_sync_blk[6] = 1'b0;
    assign proc_dep_vld_vec_0[6] = dl_detect_out ? proc_dep_vld_vec_0_reg[6] : (proc_0_data_FIFO_blk[6] | proc_0_data_PIPO_blk[6] | proc_0_start_FIFO_blk[6] | proc_0_TLF_FIFO_blk[6] | proc_0_input_sync_blk[6] | proc_0_output_sync_blk[6]);
    assign proc_0_data_FIFO_blk[7] = 1'b0 | (~kernel_pr_entry98_U0.H_write7_out_blk_n) | (~kernel_pr_entry98_U0.hyperedge_size_out7_blk_n);
    assign proc_0_data_PIPO_blk[7] = 1'b0;
    assign proc_0_start_FIFO_blk[7] = 1'b0 | (~start_for_write_back55_U0_U.if_full_n & kernel_pr_entry98_U0.ap_start & ~kernel_pr_entry98_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_write_back55_U0_U.if_read);
    assign proc_0_TLF_FIFO_blk[7] = 1'b0;
    assign proc_0_input_sync_blk[7] = 1'b0;
    assign proc_0_output_sync_blk[7] = 1'b0;
    assign proc_dep_vld_vec_0[7] = dl_detect_out ? proc_dep_vld_vec_0_reg[7] : (proc_0_data_FIFO_blk[7] | proc_0_data_PIPO_blk[7] | proc_0_start_FIFO_blk[7] | proc_0_TLF_FIFO_blk[7] | proc_0_input_sync_blk[7] | proc_0_output_sync_blk[7]);
    assign proc_0_data_FIFO_blk[8] = 1'b0 | (~kernel_pr_entry98_U0.H_write8_out_blk_n) | (~kernel_pr_entry98_U0.hyperedge_size_out8_blk_n);
    assign proc_0_data_PIPO_blk[8] = 1'b0;
    assign proc_0_start_FIFO_blk[8] = 1'b0 | (~start_for_write_back56_U0_U.if_full_n & kernel_pr_entry98_U0.ap_start & ~kernel_pr_entry98_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_write_back56_U0_U.if_read);
    assign proc_0_TLF_FIFO_blk[8] = 1'b0;
    assign proc_0_input_sync_blk[8] = 1'b0;
    assign proc_0_output_sync_blk[8] = 1'b0;
    assign proc_dep_vld_vec_0[8] = dl_detect_out ? proc_dep_vld_vec_0_reg[8] : (proc_0_data_FIFO_blk[8] | proc_0_data_PIPO_blk[8] | proc_0_start_FIFO_blk[8] | proc_0_TLF_FIFO_blk[8] | proc_0_input_sync_blk[8] | proc_0_output_sync_blk[8]);
    assign proc_0_data_FIFO_blk[9] = 1'b0 | (~kernel_pr_entry98_U0.H_write9_out_blk_n) | (~kernel_pr_entry98_U0.hyperedge_size_out9_blk_n);
    assign proc_0_data_PIPO_blk[9] = 1'b0;
    assign proc_0_start_FIFO_blk[9] = 1'b0 | (~start_for_write_back57_U0_U.if_full_n & kernel_pr_entry98_U0.ap_start & ~kernel_pr_entry98_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_write_back57_U0_U.if_read);
    assign proc_0_TLF_FIFO_blk[9] = 1'b0;
    assign proc_0_input_sync_blk[9] = 1'b0;
    assign proc_0_output_sync_blk[9] = 1'b0;
    assign proc_dep_vld_vec_0[9] = dl_detect_out ? proc_dep_vld_vec_0_reg[9] : (proc_0_data_FIFO_blk[9] | proc_0_data_PIPO_blk[9] | proc_0_start_FIFO_blk[9] | proc_0_TLF_FIFO_blk[9] | proc_0_input_sync_blk[9] | proc_0_output_sync_blk[9]);
    assign proc_0_data_FIFO_blk[10] = 1'b0 | (~kernel_pr_entry98_U0.H_write10_out_blk_n) | (~kernel_pr_entry98_U0.hyperedge_size_out10_blk_n);
    assign proc_0_data_PIPO_blk[10] = 1'b0;
    assign proc_0_start_FIFO_blk[10] = 1'b0 | (~start_for_write_back58_U0_U.if_full_n & kernel_pr_entry98_U0.ap_start & ~kernel_pr_entry98_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_write_back58_U0_U.if_read);
    assign proc_0_TLF_FIFO_blk[10] = 1'b0;
    assign proc_0_input_sync_blk[10] = 1'b0;
    assign proc_0_output_sync_blk[10] = 1'b0;
    assign proc_dep_vld_vec_0[10] = dl_detect_out ? proc_dep_vld_vec_0_reg[10] : (proc_0_data_FIFO_blk[10] | proc_0_data_PIPO_blk[10] | proc_0_start_FIFO_blk[10] | proc_0_TLF_FIFO_blk[10] | proc_0_input_sync_blk[10] | proc_0_output_sync_blk[10]);
    assign proc_0_data_FIFO_blk[11] = 1'b0 | (~kernel_pr_entry98_U0.H_write11_out_blk_n) | (~kernel_pr_entry98_U0.hyperedge_size_out11_blk_n);
    assign proc_0_data_PIPO_blk[11] = 1'b0;
    assign proc_0_start_FIFO_blk[11] = 1'b0 | (~start_for_write_back59_U0_U.if_full_n & kernel_pr_entry98_U0.ap_start & ~kernel_pr_entry98_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_write_back59_U0_U.if_read);
    assign proc_0_TLF_FIFO_blk[11] = 1'b0;
    assign proc_0_input_sync_blk[11] = 1'b0;
    assign proc_0_output_sync_blk[11] = 1'b0;
    assign proc_dep_vld_vec_0[11] = dl_detect_out ? proc_dep_vld_vec_0_reg[11] : (proc_0_data_FIFO_blk[11] | proc_0_data_PIPO_blk[11] | proc_0_start_FIFO_blk[11] | proc_0_TLF_FIFO_blk[11] | proc_0_input_sync_blk[11] | proc_0_output_sync_blk[11]);
    assign proc_0_data_FIFO_blk[12] = 1'b0 | (~kernel_pr_entry98_U0.H_write12_out_blk_n) | (~kernel_pr_entry98_U0.hyperedge_size_out12_blk_n);
    assign proc_0_data_PIPO_blk[12] = 1'b0;
    assign proc_0_start_FIFO_blk[12] = 1'b0 | (~start_for_write_back60_U0_U.if_full_n & kernel_pr_entry98_U0.ap_start & ~kernel_pr_entry98_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_write_back60_U0_U.if_read);
    assign proc_0_TLF_FIFO_blk[12] = 1'b0;
    assign proc_0_input_sync_blk[12] = 1'b0;
    assign proc_0_output_sync_blk[12] = 1'b0;
    assign proc_dep_vld_vec_0[12] = dl_detect_out ? proc_dep_vld_vec_0_reg[12] : (proc_0_data_FIFO_blk[12] | proc_0_data_PIPO_blk[12] | proc_0_start_FIFO_blk[12] | proc_0_TLF_FIFO_blk[12] | proc_0_input_sync_blk[12] | proc_0_output_sync_blk[12]);
    assign proc_0_data_FIFO_blk[13] = 1'b0 | (~kernel_pr_entry98_U0.H_write13_out_blk_n) | (~kernel_pr_entry98_U0.hyperedge_size_out13_blk_n);
    assign proc_0_data_PIPO_blk[13] = 1'b0;
    assign proc_0_start_FIFO_blk[13] = 1'b0 | (~start_for_write_back61_U0_U.if_full_n & kernel_pr_entry98_U0.ap_start & ~kernel_pr_entry98_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_write_back61_U0_U.if_read);
    assign proc_0_TLF_FIFO_blk[13] = 1'b0;
    assign proc_0_input_sync_blk[13] = 1'b0;
    assign proc_0_output_sync_blk[13] = 1'b0;
    assign proc_dep_vld_vec_0[13] = dl_detect_out ? proc_dep_vld_vec_0_reg[13] : (proc_0_data_FIFO_blk[13] | proc_0_data_PIPO_blk[13] | proc_0_start_FIFO_blk[13] | proc_0_TLF_FIFO_blk[13] | proc_0_input_sync_blk[13] | proc_0_output_sync_blk[13]);
    assign proc_0_data_FIFO_blk[14] = 1'b0 | (~kernel_pr_entry98_U0.H_write14_out_blk_n) | (~kernel_pr_entry98_U0.hyperedge_size_out14_blk_n);
    assign proc_0_data_PIPO_blk[14] = 1'b0;
    assign proc_0_start_FIFO_blk[14] = 1'b0 | (~start_for_write_back62_U0_U.if_full_n & kernel_pr_entry98_U0.ap_start & ~kernel_pr_entry98_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_write_back62_U0_U.if_read);
    assign proc_0_TLF_FIFO_blk[14] = 1'b0;
    assign proc_0_input_sync_blk[14] = 1'b0;
    assign proc_0_output_sync_blk[14] = 1'b0;
    assign proc_dep_vld_vec_0[14] = dl_detect_out ? proc_dep_vld_vec_0_reg[14] : (proc_0_data_FIFO_blk[14] | proc_0_data_PIPO_blk[14] | proc_0_start_FIFO_blk[14] | proc_0_TLF_FIFO_blk[14] | proc_0_input_sync_blk[14] | proc_0_output_sync_blk[14]);
    assign proc_0_data_FIFO_blk[15] = 1'b0 | (~kernel_pr_entry98_U0.H_write15_out_blk_n) | (~kernel_pr_entry98_U0.hyperedge_size_out15_blk_n);
    assign proc_0_data_PIPO_blk[15] = 1'b0;
    assign proc_0_start_FIFO_blk[15] = 1'b0 | (~start_for_write_back63_U0_U.if_full_n & kernel_pr_entry98_U0.ap_start & ~kernel_pr_entry98_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_write_back63_U0_U.if_read);
    assign proc_0_TLF_FIFO_blk[15] = 1'b0;
    assign proc_0_input_sync_blk[15] = 1'b0;
    assign proc_0_output_sync_blk[15] = 1'b0;
    assign proc_dep_vld_vec_0[15] = dl_detect_out ? proc_dep_vld_vec_0_reg[15] : (proc_0_data_FIFO_blk[15] | proc_0_data_PIPO_blk[15] | proc_0_start_FIFO_blk[15] | proc_0_TLF_FIFO_blk[15] | proc_0_input_sync_blk[15] | proc_0_output_sync_blk[15]);
    assign proc_0_data_FIFO_blk[16] = 1'b0 | (~kernel_pr_entry98_U0.V_read0_out_blk_n);
    assign proc_0_data_PIPO_blk[16] = 1'b0;
    assign proc_0_start_FIFO_blk[16] = 1'b0;
    assign proc_0_TLF_FIFO_blk[16] = 1'b0;
    assign proc_0_input_sync_blk[16] = 1'b0 | (ap_sync_kernel_pr_entry98_U0_ap_ready & kernel_pr_entry98_U0.ap_idle & ~ap_sync_load_value32_U0_ap_ready);
    assign proc_0_output_sync_blk[16] = 1'b0;
    assign proc_dep_vld_vec_0[16] = dl_detect_out ? proc_dep_vld_vec_0_reg[16] : (proc_0_data_FIFO_blk[16] | proc_0_data_PIPO_blk[16] | proc_0_start_FIFO_blk[16] | proc_0_TLF_FIFO_blk[16] | proc_0_input_sync_blk[16] | proc_0_output_sync_blk[16]);
    assign proc_0_data_FIFO_blk[17] = 1'b0 | (~kernel_pr_entry98_U0.V_read1_out_blk_n);
    assign proc_0_data_PIPO_blk[17] = 1'b0;
    assign proc_0_start_FIFO_blk[17] = 1'b0;
    assign proc_0_TLF_FIFO_blk[17] = 1'b0;
    assign proc_0_input_sync_blk[17] = 1'b0 | (ap_sync_kernel_pr_entry98_U0_ap_ready & kernel_pr_entry98_U0.ap_idle & ~ap_sync_load_value33_U0_ap_ready);
    assign proc_0_output_sync_blk[17] = 1'b0;
    assign proc_dep_vld_vec_0[17] = dl_detect_out ? proc_dep_vld_vec_0_reg[17] : (proc_0_data_FIFO_blk[17] | proc_0_data_PIPO_blk[17] | proc_0_start_FIFO_blk[17] | proc_0_TLF_FIFO_blk[17] | proc_0_input_sync_blk[17] | proc_0_output_sync_blk[17]);
    assign proc_0_data_FIFO_blk[18] = 1'b0 | (~kernel_pr_entry98_U0.V_read2_out_blk_n);
    assign proc_0_data_PIPO_blk[18] = 1'b0;
    assign proc_0_start_FIFO_blk[18] = 1'b0;
    assign proc_0_TLF_FIFO_blk[18] = 1'b0;
    assign proc_0_input_sync_blk[18] = 1'b0 | (ap_sync_kernel_pr_entry98_U0_ap_ready & kernel_pr_entry98_U0.ap_idle & ~ap_sync_load_value34_U0_ap_ready);
    assign proc_0_output_sync_blk[18] = 1'b0;
    assign proc_dep_vld_vec_0[18] = dl_detect_out ? proc_dep_vld_vec_0_reg[18] : (proc_0_data_FIFO_blk[18] | proc_0_data_PIPO_blk[18] | proc_0_start_FIFO_blk[18] | proc_0_TLF_FIFO_blk[18] | proc_0_input_sync_blk[18] | proc_0_output_sync_blk[18]);
    assign proc_0_data_FIFO_blk[19] = 1'b0 | (~kernel_pr_entry98_U0.V_read3_out_blk_n);
    assign proc_0_data_PIPO_blk[19] = 1'b0;
    assign proc_0_start_FIFO_blk[19] = 1'b0;
    assign proc_0_TLF_FIFO_blk[19] = 1'b0;
    assign proc_0_input_sync_blk[19] = 1'b0 | (ap_sync_kernel_pr_entry98_U0_ap_ready & kernel_pr_entry98_U0.ap_idle & ~ap_sync_load_value35_U0_ap_ready);
    assign proc_0_output_sync_blk[19] = 1'b0;
    assign proc_dep_vld_vec_0[19] = dl_detect_out ? proc_dep_vld_vec_0_reg[19] : (proc_0_data_FIFO_blk[19] | proc_0_data_PIPO_blk[19] | proc_0_start_FIFO_blk[19] | proc_0_TLF_FIFO_blk[19] | proc_0_input_sync_blk[19] | proc_0_output_sync_blk[19]);
    assign proc_0_data_FIFO_blk[20] = 1'b0 | (~kernel_pr_entry98_U0.V_read4_out_blk_n);
    assign proc_0_data_PIPO_blk[20] = 1'b0;
    assign proc_0_start_FIFO_blk[20] = 1'b0;
    assign proc_0_TLF_FIFO_blk[20] = 1'b0;
    assign proc_0_input_sync_blk[20] = 1'b0 | (ap_sync_kernel_pr_entry98_U0_ap_ready & kernel_pr_entry98_U0.ap_idle & ~ap_sync_load_value36_U0_ap_ready);
    assign proc_0_output_sync_blk[20] = 1'b0;
    assign proc_dep_vld_vec_0[20] = dl_detect_out ? proc_dep_vld_vec_0_reg[20] : (proc_0_data_FIFO_blk[20] | proc_0_data_PIPO_blk[20] | proc_0_start_FIFO_blk[20] | proc_0_TLF_FIFO_blk[20] | proc_0_input_sync_blk[20] | proc_0_output_sync_blk[20]);
    assign proc_0_data_FIFO_blk[21] = 1'b0 | (~kernel_pr_entry98_U0.V_read5_out_blk_n);
    assign proc_0_data_PIPO_blk[21] = 1'b0;
    assign proc_0_start_FIFO_blk[21] = 1'b0;
    assign proc_0_TLF_FIFO_blk[21] = 1'b0;
    assign proc_0_input_sync_blk[21] = 1'b0 | (ap_sync_kernel_pr_entry98_U0_ap_ready & kernel_pr_entry98_U0.ap_idle & ~ap_sync_load_value37_U0_ap_ready);
    assign proc_0_output_sync_blk[21] = 1'b0;
    assign proc_dep_vld_vec_0[21] = dl_detect_out ? proc_dep_vld_vec_0_reg[21] : (proc_0_data_FIFO_blk[21] | proc_0_data_PIPO_blk[21] | proc_0_start_FIFO_blk[21] | proc_0_TLF_FIFO_blk[21] | proc_0_input_sync_blk[21] | proc_0_output_sync_blk[21]);
    assign proc_0_data_FIFO_blk[22] = 1'b0 | (~kernel_pr_entry98_U0.V_read6_out_blk_n);
    assign proc_0_data_PIPO_blk[22] = 1'b0;
    assign proc_0_start_FIFO_blk[22] = 1'b0;
    assign proc_0_TLF_FIFO_blk[22] = 1'b0;
    assign proc_0_input_sync_blk[22] = 1'b0 | (ap_sync_kernel_pr_entry98_U0_ap_ready & kernel_pr_entry98_U0.ap_idle & ~ap_sync_load_value38_U0_ap_ready);
    assign proc_0_output_sync_blk[22] = 1'b0;
    assign proc_dep_vld_vec_0[22] = dl_detect_out ? proc_dep_vld_vec_0_reg[22] : (proc_0_data_FIFO_blk[22] | proc_0_data_PIPO_blk[22] | proc_0_start_FIFO_blk[22] | proc_0_TLF_FIFO_blk[22] | proc_0_input_sync_blk[22] | proc_0_output_sync_blk[22]);
    assign proc_0_data_FIFO_blk[23] = 1'b0 | (~kernel_pr_entry98_U0.V_read7_out_blk_n);
    assign proc_0_data_PIPO_blk[23] = 1'b0;
    assign proc_0_start_FIFO_blk[23] = 1'b0;
    assign proc_0_TLF_FIFO_blk[23] = 1'b0;
    assign proc_0_input_sync_blk[23] = 1'b0 | (ap_sync_kernel_pr_entry98_U0_ap_ready & kernel_pr_entry98_U0.ap_idle & ~ap_sync_load_value39_U0_ap_ready);
    assign proc_0_output_sync_blk[23] = 1'b0;
    assign proc_dep_vld_vec_0[23] = dl_detect_out ? proc_dep_vld_vec_0_reg[23] : (proc_0_data_FIFO_blk[23] | proc_0_data_PIPO_blk[23] | proc_0_start_FIFO_blk[23] | proc_0_TLF_FIFO_blk[23] | proc_0_input_sync_blk[23] | proc_0_output_sync_blk[23]);
    assign proc_0_data_FIFO_blk[24] = 1'b0 | (~kernel_pr_entry98_U0.V_read8_out_blk_n);
    assign proc_0_data_PIPO_blk[24] = 1'b0;
    assign proc_0_start_FIFO_blk[24] = 1'b0;
    assign proc_0_TLF_FIFO_blk[24] = 1'b0;
    assign proc_0_input_sync_blk[24] = 1'b0 | (ap_sync_kernel_pr_entry98_U0_ap_ready & kernel_pr_entry98_U0.ap_idle & ~ap_sync_load_value40_U0_ap_ready);
    assign proc_0_output_sync_blk[24] = 1'b0;
    assign proc_dep_vld_vec_0[24] = dl_detect_out ? proc_dep_vld_vec_0_reg[24] : (proc_0_data_FIFO_blk[24] | proc_0_data_PIPO_blk[24] | proc_0_start_FIFO_blk[24] | proc_0_TLF_FIFO_blk[24] | proc_0_input_sync_blk[24] | proc_0_output_sync_blk[24]);
    assign proc_0_data_FIFO_blk[25] = 1'b0 | (~kernel_pr_entry98_U0.V_read9_out_blk_n);
    assign proc_0_data_PIPO_blk[25] = 1'b0;
    assign proc_0_start_FIFO_blk[25] = 1'b0;
    assign proc_0_TLF_FIFO_blk[25] = 1'b0;
    assign proc_0_input_sync_blk[25] = 1'b0 | (ap_sync_kernel_pr_entry98_U0_ap_ready & kernel_pr_entry98_U0.ap_idle & ~ap_sync_load_value41_U0_ap_ready);
    assign proc_0_output_sync_blk[25] = 1'b0;
    assign proc_dep_vld_vec_0[25] = dl_detect_out ? proc_dep_vld_vec_0_reg[25] : (proc_0_data_FIFO_blk[25] | proc_0_data_PIPO_blk[25] | proc_0_start_FIFO_blk[25] | proc_0_TLF_FIFO_blk[25] | proc_0_input_sync_blk[25] | proc_0_output_sync_blk[25]);
    assign proc_0_data_FIFO_blk[26] = 1'b0 | (~kernel_pr_entry98_U0.V_read10_out_blk_n);
    assign proc_0_data_PIPO_blk[26] = 1'b0;
    assign proc_0_start_FIFO_blk[26] = 1'b0;
    assign proc_0_TLF_FIFO_blk[26] = 1'b0;
    assign proc_0_input_sync_blk[26] = 1'b0 | (ap_sync_kernel_pr_entry98_U0_ap_ready & kernel_pr_entry98_U0.ap_idle & ~ap_sync_load_value42_U0_ap_ready);
    assign proc_0_output_sync_blk[26] = 1'b0;
    assign proc_dep_vld_vec_0[26] = dl_detect_out ? proc_dep_vld_vec_0_reg[26] : (proc_0_data_FIFO_blk[26] | proc_0_data_PIPO_blk[26] | proc_0_start_FIFO_blk[26] | proc_0_TLF_FIFO_blk[26] | proc_0_input_sync_blk[26] | proc_0_output_sync_blk[26]);
    assign proc_0_data_FIFO_blk[27] = 1'b0 | (~kernel_pr_entry98_U0.V_read11_out_blk_n);
    assign proc_0_data_PIPO_blk[27] = 1'b0;
    assign proc_0_start_FIFO_blk[27] = 1'b0;
    assign proc_0_TLF_FIFO_blk[27] = 1'b0;
    assign proc_0_input_sync_blk[27] = 1'b0 | (ap_sync_kernel_pr_entry98_U0_ap_ready & kernel_pr_entry98_U0.ap_idle & ~ap_sync_load_value43_U0_ap_ready);
    assign proc_0_output_sync_blk[27] = 1'b0;
    assign proc_dep_vld_vec_0[27] = dl_detect_out ? proc_dep_vld_vec_0_reg[27] : (proc_0_data_FIFO_blk[27] | proc_0_data_PIPO_blk[27] | proc_0_start_FIFO_blk[27] | proc_0_TLF_FIFO_blk[27] | proc_0_input_sync_blk[27] | proc_0_output_sync_blk[27]);
    assign proc_0_data_FIFO_blk[28] = 1'b0 | (~kernel_pr_entry98_U0.V_read12_out_blk_n);
    assign proc_0_data_PIPO_blk[28] = 1'b0;
    assign proc_0_start_FIFO_blk[28] = 1'b0;
    assign proc_0_TLF_FIFO_blk[28] = 1'b0;
    assign proc_0_input_sync_blk[28] = 1'b0 | (ap_sync_kernel_pr_entry98_U0_ap_ready & kernel_pr_entry98_U0.ap_idle & ~ap_sync_load_value44_U0_ap_ready);
    assign proc_0_output_sync_blk[28] = 1'b0;
    assign proc_dep_vld_vec_0[28] = dl_detect_out ? proc_dep_vld_vec_0_reg[28] : (proc_0_data_FIFO_blk[28] | proc_0_data_PIPO_blk[28] | proc_0_start_FIFO_blk[28] | proc_0_TLF_FIFO_blk[28] | proc_0_input_sync_blk[28] | proc_0_output_sync_blk[28]);
    assign proc_0_data_FIFO_blk[29] = 1'b0 | (~kernel_pr_entry98_U0.V_read13_out_blk_n);
    assign proc_0_data_PIPO_blk[29] = 1'b0;
    assign proc_0_start_FIFO_blk[29] = 1'b0;
    assign proc_0_TLF_FIFO_blk[29] = 1'b0;
    assign proc_0_input_sync_blk[29] = 1'b0 | (ap_sync_kernel_pr_entry98_U0_ap_ready & kernel_pr_entry98_U0.ap_idle & ~ap_sync_load_value45_U0_ap_ready);
    assign proc_0_output_sync_blk[29] = 1'b0;
    assign proc_dep_vld_vec_0[29] = dl_detect_out ? proc_dep_vld_vec_0_reg[29] : (proc_0_data_FIFO_blk[29] | proc_0_data_PIPO_blk[29] | proc_0_start_FIFO_blk[29] | proc_0_TLF_FIFO_blk[29] | proc_0_input_sync_blk[29] | proc_0_output_sync_blk[29]);
    assign proc_0_data_FIFO_blk[30] = 1'b0 | (~kernel_pr_entry98_U0.V_read14_out_blk_n);
    assign proc_0_data_PIPO_blk[30] = 1'b0;
    assign proc_0_start_FIFO_blk[30] = 1'b0;
    assign proc_0_TLF_FIFO_blk[30] = 1'b0;
    assign proc_0_input_sync_blk[30] = 1'b0 | (ap_sync_kernel_pr_entry98_U0_ap_ready & kernel_pr_entry98_U0.ap_idle & ~ap_sync_load_value46_U0_ap_ready);
    assign proc_0_output_sync_blk[30] = 1'b0;
    assign proc_dep_vld_vec_0[30] = dl_detect_out ? proc_dep_vld_vec_0_reg[30] : (proc_0_data_FIFO_blk[30] | proc_0_data_PIPO_blk[30] | proc_0_start_FIFO_blk[30] | proc_0_TLF_FIFO_blk[30] | proc_0_input_sync_blk[30] | proc_0_output_sync_blk[30]);
    assign proc_0_data_FIFO_blk[31] = 1'b0 | (~kernel_pr_entry98_U0.V_read15_out_blk_n);
    assign proc_0_data_PIPO_blk[31] = 1'b0;
    assign proc_0_start_FIFO_blk[31] = 1'b0;
    assign proc_0_TLF_FIFO_blk[31] = 1'b0;
    assign proc_0_input_sync_blk[31] = 1'b0 | (ap_sync_kernel_pr_entry98_U0_ap_ready & kernel_pr_entry98_U0.ap_idle & ~ap_sync_load_value47_U0_ap_ready);
    assign proc_0_output_sync_blk[31] = 1'b0;
    assign proc_dep_vld_vec_0[31] = dl_detect_out ? proc_dep_vld_vec_0_reg[31] : (proc_0_data_FIFO_blk[31] | proc_0_data_PIPO_blk[31] | proc_0_start_FIFO_blk[31] | proc_0_TLF_FIFO_blk[31] | proc_0_input_sync_blk[31] | proc_0_output_sync_blk[31]);
    assign proc_0_data_FIFO_blk[32] = 1'b0 | (~kernel_pr_entry98_U0.hv_bipedge_dram0_out_blk_n) | (~kernel_pr_entry98_U0.bipedge_size_out_blk_n);
    assign proc_0_data_PIPO_blk[32] = 1'b0;
    assign proc_0_start_FIFO_blk[32] = 1'b0;
    assign proc_0_TLF_FIFO_blk[32] = 1'b0;
    assign proc_0_input_sync_blk[32] = 1'b0 | (ap_sync_kernel_pr_entry98_U0_ap_ready & kernel_pr_entry98_U0.ap_idle & ~ap_sync_load_bipedge30_U0_ap_ready);
    assign proc_0_output_sync_blk[32] = 1'b0;
    assign proc_dep_vld_vec_0[32] = dl_detect_out ? proc_dep_vld_vec_0_reg[32] : (proc_0_data_FIFO_blk[32] | proc_0_data_PIPO_blk[32] | proc_0_start_FIFO_blk[32] | proc_0_TLF_FIFO_blk[32] | proc_0_input_sync_blk[32] | proc_0_output_sync_blk[32]);
    assign proc_0_data_FIFO_blk[33] = 1'b0 | (~kernel_pr_entry98_U0.hv_bipedge_dram1_out_blk_n) | (~kernel_pr_entry98_U0.bipedge_size_out16_blk_n);
    assign proc_0_data_PIPO_blk[33] = 1'b0;
    assign proc_0_start_FIFO_blk[33] = 1'b0;
    assign proc_0_TLF_FIFO_blk[33] = 1'b0;
    assign proc_0_input_sync_blk[33] = 1'b0 | (ap_sync_kernel_pr_entry98_U0_ap_ready & kernel_pr_entry98_U0.ap_idle & ~ap_sync_load_bipedge31_U0_ap_ready);
    assign proc_0_output_sync_blk[33] = 1'b0;
    assign proc_dep_vld_vec_0[33] = dl_detect_out ? proc_dep_vld_vec_0_reg[33] : (proc_0_data_FIFO_blk[33] | proc_0_data_PIPO_blk[33] | proc_0_start_FIFO_blk[33] | proc_0_TLF_FIFO_blk[33] | proc_0_input_sync_blk[33] | proc_0_output_sync_blk[33]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_0_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_0_reg <= proc_dep_vld_vec_0;
        end
    end
    assign in_chan_dep_vld_vec_0[0] = dep_chan_vld_1_0;
    assign in_chan_dep_data_vec_0[34 : 0] = dep_chan_data_1_0;
    assign token_in_vec_0[0] = token_1_0;
    assign in_chan_dep_vld_vec_0[1] = dep_chan_vld_2_0;
    assign in_chan_dep_data_vec_0[69 : 35] = dep_chan_data_2_0;
    assign token_in_vec_0[1] = token_2_0;
    assign in_chan_dep_vld_vec_0[2] = dep_chan_vld_3_0;
    assign in_chan_dep_data_vec_0[104 : 70] = dep_chan_data_3_0;
    assign token_in_vec_0[2] = token_3_0;
    assign in_chan_dep_vld_vec_0[3] = dep_chan_vld_4_0;
    assign in_chan_dep_data_vec_0[139 : 105] = dep_chan_data_4_0;
    assign token_in_vec_0[3] = token_4_0;
    assign in_chan_dep_vld_vec_0[4] = dep_chan_vld_5_0;
    assign in_chan_dep_data_vec_0[174 : 140] = dep_chan_data_5_0;
    assign token_in_vec_0[4] = token_5_0;
    assign in_chan_dep_vld_vec_0[5] = dep_chan_vld_6_0;
    assign in_chan_dep_data_vec_0[209 : 175] = dep_chan_data_6_0;
    assign token_in_vec_0[5] = token_6_0;
    assign in_chan_dep_vld_vec_0[6] = dep_chan_vld_7_0;
    assign in_chan_dep_data_vec_0[244 : 210] = dep_chan_data_7_0;
    assign token_in_vec_0[6] = token_7_0;
    assign in_chan_dep_vld_vec_0[7] = dep_chan_vld_8_0;
    assign in_chan_dep_data_vec_0[279 : 245] = dep_chan_data_8_0;
    assign token_in_vec_0[7] = token_8_0;
    assign in_chan_dep_vld_vec_0[8] = dep_chan_vld_9_0;
    assign in_chan_dep_data_vec_0[314 : 280] = dep_chan_data_9_0;
    assign token_in_vec_0[8] = token_9_0;
    assign in_chan_dep_vld_vec_0[9] = dep_chan_vld_10_0;
    assign in_chan_dep_data_vec_0[349 : 315] = dep_chan_data_10_0;
    assign token_in_vec_0[9] = token_10_0;
    assign in_chan_dep_vld_vec_0[10] = dep_chan_vld_11_0;
    assign in_chan_dep_data_vec_0[384 : 350] = dep_chan_data_11_0;
    assign token_in_vec_0[10] = token_11_0;
    assign in_chan_dep_vld_vec_0[11] = dep_chan_vld_12_0;
    assign in_chan_dep_data_vec_0[419 : 385] = dep_chan_data_12_0;
    assign token_in_vec_0[11] = token_12_0;
    assign in_chan_dep_vld_vec_0[12] = dep_chan_vld_13_0;
    assign in_chan_dep_data_vec_0[454 : 420] = dep_chan_data_13_0;
    assign token_in_vec_0[12] = token_13_0;
    assign in_chan_dep_vld_vec_0[13] = dep_chan_vld_14_0;
    assign in_chan_dep_data_vec_0[489 : 455] = dep_chan_data_14_0;
    assign token_in_vec_0[13] = token_14_0;
    assign in_chan_dep_vld_vec_0[14] = dep_chan_vld_15_0;
    assign in_chan_dep_data_vec_0[524 : 490] = dep_chan_data_15_0;
    assign token_in_vec_0[14] = token_15_0;
    assign in_chan_dep_vld_vec_0[15] = dep_chan_vld_16_0;
    assign in_chan_dep_data_vec_0[559 : 525] = dep_chan_data_16_0;
    assign token_in_vec_0[15] = token_16_0;
    assign in_chan_dep_vld_vec_0[16] = dep_chan_vld_17_0;
    assign in_chan_dep_data_vec_0[594 : 560] = dep_chan_data_17_0;
    assign token_in_vec_0[16] = token_17_0;
    assign in_chan_dep_vld_vec_0[17] = dep_chan_vld_18_0;
    assign in_chan_dep_data_vec_0[629 : 595] = dep_chan_data_18_0;
    assign token_in_vec_0[17] = token_18_0;
    assign in_chan_dep_vld_vec_0[18] = dep_chan_vld_19_0;
    assign in_chan_dep_data_vec_0[664 : 630] = dep_chan_data_19_0;
    assign token_in_vec_0[18] = token_19_0;
    assign in_chan_dep_vld_vec_0[19] = dep_chan_vld_20_0;
    assign in_chan_dep_data_vec_0[699 : 665] = dep_chan_data_20_0;
    assign token_in_vec_0[19] = token_20_0;
    assign in_chan_dep_vld_vec_0[20] = dep_chan_vld_21_0;
    assign in_chan_dep_data_vec_0[734 : 700] = dep_chan_data_21_0;
    assign token_in_vec_0[20] = token_21_0;
    assign in_chan_dep_vld_vec_0[21] = dep_chan_vld_22_0;
    assign in_chan_dep_data_vec_0[769 : 735] = dep_chan_data_22_0;
    assign token_in_vec_0[21] = token_22_0;
    assign in_chan_dep_vld_vec_0[22] = dep_chan_vld_23_0;
    assign in_chan_dep_data_vec_0[804 : 770] = dep_chan_data_23_0;
    assign token_in_vec_0[22] = token_23_0;
    assign in_chan_dep_vld_vec_0[23] = dep_chan_vld_24_0;
    assign in_chan_dep_data_vec_0[839 : 805] = dep_chan_data_24_0;
    assign token_in_vec_0[23] = token_24_0;
    assign in_chan_dep_vld_vec_0[24] = dep_chan_vld_25_0;
    assign in_chan_dep_data_vec_0[874 : 840] = dep_chan_data_25_0;
    assign token_in_vec_0[24] = token_25_0;
    assign in_chan_dep_vld_vec_0[25] = dep_chan_vld_26_0;
    assign in_chan_dep_data_vec_0[909 : 875] = dep_chan_data_26_0;
    assign token_in_vec_0[25] = token_26_0;
    assign in_chan_dep_vld_vec_0[26] = dep_chan_vld_27_0;
    assign in_chan_dep_data_vec_0[944 : 910] = dep_chan_data_27_0;
    assign token_in_vec_0[26] = token_27_0;
    assign in_chan_dep_vld_vec_0[27] = dep_chan_vld_28_0;
    assign in_chan_dep_data_vec_0[979 : 945] = dep_chan_data_28_0;
    assign token_in_vec_0[27] = token_28_0;
    assign in_chan_dep_vld_vec_0[28] = dep_chan_vld_29_0;
    assign in_chan_dep_data_vec_0[1014 : 980] = dep_chan_data_29_0;
    assign token_in_vec_0[28] = token_29_0;
    assign in_chan_dep_vld_vec_0[29] = dep_chan_vld_30_0;
    assign in_chan_dep_data_vec_0[1049 : 1015] = dep_chan_data_30_0;
    assign token_in_vec_0[29] = token_30_0;
    assign in_chan_dep_vld_vec_0[30] = dep_chan_vld_31_0;
    assign in_chan_dep_data_vec_0[1084 : 1050] = dep_chan_data_31_0;
    assign token_in_vec_0[30] = token_31_0;
    assign in_chan_dep_vld_vec_0[31] = dep_chan_vld_32_0;
    assign in_chan_dep_data_vec_0[1119 : 1085] = dep_chan_data_32_0;
    assign token_in_vec_0[31] = token_32_0;
    assign in_chan_dep_vld_vec_0[32] = dep_chan_vld_33_0;
    assign in_chan_dep_data_vec_0[1154 : 1120] = dep_chan_data_33_0;
    assign token_in_vec_0[32] = token_33_0;
    assign in_chan_dep_vld_vec_0[33] = dep_chan_vld_34_0;
    assign in_chan_dep_data_vec_0[1189 : 1155] = dep_chan_data_34_0;
    assign token_in_vec_0[33] = token_34_0;
    assign dep_chan_vld_0_19 = out_chan_dep_vld_vec_0[0];
    assign dep_chan_data_0_19 = out_chan_dep_data_0;
    assign token_0_19 = token_out_vec_0[0];
    assign dep_chan_vld_0_20 = out_chan_dep_vld_vec_0[1];
    assign dep_chan_data_0_20 = out_chan_dep_data_0;
    assign token_0_20 = token_out_vec_0[1];
    assign dep_chan_vld_0_21 = out_chan_dep_vld_vec_0[2];
    assign dep_chan_data_0_21 = out_chan_dep_data_0;
    assign token_0_21 = token_out_vec_0[2];
    assign dep_chan_vld_0_22 = out_chan_dep_vld_vec_0[3];
    assign dep_chan_data_0_22 = out_chan_dep_data_0;
    assign token_0_22 = token_out_vec_0[3];
    assign dep_chan_vld_0_23 = out_chan_dep_vld_vec_0[4];
    assign dep_chan_data_0_23 = out_chan_dep_data_0;
    assign token_0_23 = token_out_vec_0[4];
    assign dep_chan_vld_0_24 = out_chan_dep_vld_vec_0[5];
    assign dep_chan_data_0_24 = out_chan_dep_data_0;
    assign token_0_24 = token_out_vec_0[5];
    assign dep_chan_vld_0_25 = out_chan_dep_vld_vec_0[6];
    assign dep_chan_data_0_25 = out_chan_dep_data_0;
    assign token_0_25 = token_out_vec_0[6];
    assign dep_chan_vld_0_26 = out_chan_dep_vld_vec_0[7];
    assign dep_chan_data_0_26 = out_chan_dep_data_0;
    assign token_0_26 = token_out_vec_0[7];
    assign dep_chan_vld_0_27 = out_chan_dep_vld_vec_0[8];
    assign dep_chan_data_0_27 = out_chan_dep_data_0;
    assign token_0_27 = token_out_vec_0[8];
    assign dep_chan_vld_0_28 = out_chan_dep_vld_vec_0[9];
    assign dep_chan_data_0_28 = out_chan_dep_data_0;
    assign token_0_28 = token_out_vec_0[9];
    assign dep_chan_vld_0_29 = out_chan_dep_vld_vec_0[10];
    assign dep_chan_data_0_29 = out_chan_dep_data_0;
    assign token_0_29 = token_out_vec_0[10];
    assign dep_chan_vld_0_30 = out_chan_dep_vld_vec_0[11];
    assign dep_chan_data_0_30 = out_chan_dep_data_0;
    assign token_0_30 = token_out_vec_0[11];
    assign dep_chan_vld_0_31 = out_chan_dep_vld_vec_0[12];
    assign dep_chan_data_0_31 = out_chan_dep_data_0;
    assign token_0_31 = token_out_vec_0[12];
    assign dep_chan_vld_0_32 = out_chan_dep_vld_vec_0[13];
    assign dep_chan_data_0_32 = out_chan_dep_data_0;
    assign token_0_32 = token_out_vec_0[13];
    assign dep_chan_vld_0_33 = out_chan_dep_vld_vec_0[14];
    assign dep_chan_data_0_33 = out_chan_dep_data_0;
    assign token_0_33 = token_out_vec_0[14];
    assign dep_chan_vld_0_34 = out_chan_dep_vld_vec_0[15];
    assign dep_chan_data_0_34 = out_chan_dep_data_0;
    assign token_0_34 = token_out_vec_0[15];
    assign dep_chan_vld_0_3 = out_chan_dep_vld_vec_0[16];
    assign dep_chan_data_0_3 = out_chan_dep_data_0;
    assign token_0_3 = token_out_vec_0[16];
    assign dep_chan_vld_0_4 = out_chan_dep_vld_vec_0[17];
    assign dep_chan_data_0_4 = out_chan_dep_data_0;
    assign token_0_4 = token_out_vec_0[17];
    assign dep_chan_vld_0_5 = out_chan_dep_vld_vec_0[18];
    assign dep_chan_data_0_5 = out_chan_dep_data_0;
    assign token_0_5 = token_out_vec_0[18];
    assign dep_chan_vld_0_6 = out_chan_dep_vld_vec_0[19];
    assign dep_chan_data_0_6 = out_chan_dep_data_0;
    assign token_0_6 = token_out_vec_0[19];
    assign dep_chan_vld_0_7 = out_chan_dep_vld_vec_0[20];
    assign dep_chan_data_0_7 = out_chan_dep_data_0;
    assign token_0_7 = token_out_vec_0[20];
    assign dep_chan_vld_0_8 = out_chan_dep_vld_vec_0[21];
    assign dep_chan_data_0_8 = out_chan_dep_data_0;
    assign token_0_8 = token_out_vec_0[21];
    assign dep_chan_vld_0_9 = out_chan_dep_vld_vec_0[22];
    assign dep_chan_data_0_9 = out_chan_dep_data_0;
    assign token_0_9 = token_out_vec_0[22];
    assign dep_chan_vld_0_10 = out_chan_dep_vld_vec_0[23];
    assign dep_chan_data_0_10 = out_chan_dep_data_0;
    assign token_0_10 = token_out_vec_0[23];
    assign dep_chan_vld_0_11 = out_chan_dep_vld_vec_0[24];
    assign dep_chan_data_0_11 = out_chan_dep_data_0;
    assign token_0_11 = token_out_vec_0[24];
    assign dep_chan_vld_0_12 = out_chan_dep_vld_vec_0[25];
    assign dep_chan_data_0_12 = out_chan_dep_data_0;
    assign token_0_12 = token_out_vec_0[25];
    assign dep_chan_vld_0_13 = out_chan_dep_vld_vec_0[26];
    assign dep_chan_data_0_13 = out_chan_dep_data_0;
    assign token_0_13 = token_out_vec_0[26];
    assign dep_chan_vld_0_14 = out_chan_dep_vld_vec_0[27];
    assign dep_chan_data_0_14 = out_chan_dep_data_0;
    assign token_0_14 = token_out_vec_0[27];
    assign dep_chan_vld_0_15 = out_chan_dep_vld_vec_0[28];
    assign dep_chan_data_0_15 = out_chan_dep_data_0;
    assign token_0_15 = token_out_vec_0[28];
    assign dep_chan_vld_0_16 = out_chan_dep_vld_vec_0[29];
    assign dep_chan_data_0_16 = out_chan_dep_data_0;
    assign token_0_16 = token_out_vec_0[29];
    assign dep_chan_vld_0_17 = out_chan_dep_vld_vec_0[30];
    assign dep_chan_data_0_17 = out_chan_dep_data_0;
    assign token_0_17 = token_out_vec_0[30];
    assign dep_chan_vld_0_18 = out_chan_dep_vld_vec_0[31];
    assign dep_chan_data_0_18 = out_chan_dep_data_0;
    assign token_0_18 = token_out_vec_0[31];
    assign dep_chan_vld_0_1 = out_chan_dep_vld_vec_0[32];
    assign dep_chan_data_0_1 = out_chan_dep_data_0;
    assign token_0_1 = token_out_vec_0[32];
    assign dep_chan_vld_0_2 = out_chan_dep_vld_vec_0[33];
    assign dep_chan_data_0_2 = out_chan_dep_data_0;
    assign token_0_2 = token_out_vec_0[33];

    // Process: load_bipedge30_U0
    kernel_pr_hls_deadlock_detect_unit #(35, 1, 18, 18) kernel_pr_hls_deadlock_detect_unit_1 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_1),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_1),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_1),
        .token_in_vec(token_in_vec_1),
        .dl_detect_in(dl_detect_out),
        .origin(origin[1]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_1),
        .out_chan_dep_data(out_chan_dep_data_1),
        .token_out_vec(token_out_vec_1),
        .dl_detect_out(dl_in_vec[1]));

    assign proc_1_data_FIFO_blk[0] = 1'b0 | (~load_bipedge30_U0.bipedge_blk_n) | (~load_bipedge30_U0.bipedge_size_blk_n);
    assign proc_1_data_PIPO_blk[0] = 1'b0;
    assign proc_1_start_FIFO_blk[0] = 1'b0;
    assign proc_1_TLF_FIFO_blk[0] = 1'b0;
    assign proc_1_input_sync_blk[0] = 1'b0 | (ap_sync_load_bipedge30_U0_ap_ready & load_bipedge30_U0.ap_idle & ~ap_sync_kernel_pr_entry98_U0_ap_ready);
    assign proc_1_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_1[0] = dl_detect_out ? proc_dep_vld_vec_1_reg[0] : (proc_1_data_FIFO_blk[0] | proc_1_data_PIPO_blk[0] | proc_1_start_FIFO_blk[0] | proc_1_TLF_FIFO_blk[0] | proc_1_input_sync_blk[0] | proc_1_output_sync_blk[0]);
    assign proc_1_data_FIFO_blk[1] = 1'b0 | (~load_bipedge30_U0.bipedge_stream_blk_n) | (~load_bipedge30_U0.bipedge_size_out_blk_n);
    assign proc_1_data_PIPO_blk[1] = 1'b0;
    assign proc_1_start_FIFO_blk[1] = 1'b0;
    assign proc_1_TLF_FIFO_blk[1] = 1'b0;
    assign proc_1_input_sync_blk[1] = 1'b0 | (ap_sync_load_bipedge30_U0_ap_ready & load_bipedge30_U0.ap_idle & ~ap_sync_load_value32_U0_ap_ready);
    assign proc_1_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_1[1] = dl_detect_out ? proc_dep_vld_vec_1_reg[1] : (proc_1_data_FIFO_blk[1] | proc_1_data_PIPO_blk[1] | proc_1_start_FIFO_blk[1] | proc_1_TLF_FIFO_blk[1] | proc_1_input_sync_blk[1] | proc_1_output_sync_blk[1]);
    assign proc_1_data_FIFO_blk[2] = 1'b0 | (~load_bipedge30_U0.bipedge_stream1_blk_n) | (~load_bipedge30_U0.bipedge_size_out1_blk_n);
    assign proc_1_data_PIPO_blk[2] = 1'b0;
    assign proc_1_start_FIFO_blk[2] = 1'b0;
    assign proc_1_TLF_FIFO_blk[2] = 1'b0;
    assign proc_1_input_sync_blk[2] = 1'b0 | (ap_sync_load_bipedge30_U0_ap_ready & load_bipedge30_U0.ap_idle & ~ap_sync_load_value33_U0_ap_ready);
    assign proc_1_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_1[2] = dl_detect_out ? proc_dep_vld_vec_1_reg[2] : (proc_1_data_FIFO_blk[2] | proc_1_data_PIPO_blk[2] | proc_1_start_FIFO_blk[2] | proc_1_TLF_FIFO_blk[2] | proc_1_input_sync_blk[2] | proc_1_output_sync_blk[2]);
    assign proc_1_data_FIFO_blk[3] = 1'b0 | (~load_bipedge30_U0.bipedge_stream2_blk_n) | (~load_bipedge30_U0.bipedge_size_out2_blk_n);
    assign proc_1_data_PIPO_blk[3] = 1'b0;
    assign proc_1_start_FIFO_blk[3] = 1'b0;
    assign proc_1_TLF_FIFO_blk[3] = 1'b0;
    assign proc_1_input_sync_blk[3] = 1'b0 | (ap_sync_load_bipedge30_U0_ap_ready & load_bipedge30_U0.ap_idle & ~ap_sync_load_value34_U0_ap_ready);
    assign proc_1_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_1[3] = dl_detect_out ? proc_dep_vld_vec_1_reg[3] : (proc_1_data_FIFO_blk[3] | proc_1_data_PIPO_blk[3] | proc_1_start_FIFO_blk[3] | proc_1_TLF_FIFO_blk[3] | proc_1_input_sync_blk[3] | proc_1_output_sync_blk[3]);
    assign proc_1_data_FIFO_blk[4] = 1'b0 | (~load_bipedge30_U0.bipedge_stream3_blk_n) | (~load_bipedge30_U0.bipedge_size_out3_blk_n);
    assign proc_1_data_PIPO_blk[4] = 1'b0;
    assign proc_1_start_FIFO_blk[4] = 1'b0;
    assign proc_1_TLF_FIFO_blk[4] = 1'b0;
    assign proc_1_input_sync_blk[4] = 1'b0 | (ap_sync_load_bipedge30_U0_ap_ready & load_bipedge30_U0.ap_idle & ~ap_sync_load_value35_U0_ap_ready);
    assign proc_1_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_1[4] = dl_detect_out ? proc_dep_vld_vec_1_reg[4] : (proc_1_data_FIFO_blk[4] | proc_1_data_PIPO_blk[4] | proc_1_start_FIFO_blk[4] | proc_1_TLF_FIFO_blk[4] | proc_1_input_sync_blk[4] | proc_1_output_sync_blk[4]);
    assign proc_1_data_FIFO_blk[5] = 1'b0 | (~load_bipedge30_U0.bipedge_stream4_blk_n) | (~load_bipedge30_U0.bipedge_size_out4_blk_n);
    assign proc_1_data_PIPO_blk[5] = 1'b0;
    assign proc_1_start_FIFO_blk[5] = 1'b0;
    assign proc_1_TLF_FIFO_blk[5] = 1'b0;
    assign proc_1_input_sync_blk[5] = 1'b0 | (ap_sync_load_bipedge30_U0_ap_ready & load_bipedge30_U0.ap_idle & ~ap_sync_load_value36_U0_ap_ready);
    assign proc_1_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_1[5] = dl_detect_out ? proc_dep_vld_vec_1_reg[5] : (proc_1_data_FIFO_blk[5] | proc_1_data_PIPO_blk[5] | proc_1_start_FIFO_blk[5] | proc_1_TLF_FIFO_blk[5] | proc_1_input_sync_blk[5] | proc_1_output_sync_blk[5]);
    assign proc_1_data_FIFO_blk[6] = 1'b0 | (~load_bipedge30_U0.bipedge_stream5_blk_n) | (~load_bipedge30_U0.bipedge_size_out5_blk_n);
    assign proc_1_data_PIPO_blk[6] = 1'b0;
    assign proc_1_start_FIFO_blk[6] = 1'b0;
    assign proc_1_TLF_FIFO_blk[6] = 1'b0;
    assign proc_1_input_sync_blk[6] = 1'b0 | (ap_sync_load_bipedge30_U0_ap_ready & load_bipedge30_U0.ap_idle & ~ap_sync_load_value37_U0_ap_ready);
    assign proc_1_output_sync_blk[6] = 1'b0;
    assign proc_dep_vld_vec_1[6] = dl_detect_out ? proc_dep_vld_vec_1_reg[6] : (proc_1_data_FIFO_blk[6] | proc_1_data_PIPO_blk[6] | proc_1_start_FIFO_blk[6] | proc_1_TLF_FIFO_blk[6] | proc_1_input_sync_blk[6] | proc_1_output_sync_blk[6]);
    assign proc_1_data_FIFO_blk[7] = 1'b0 | (~load_bipedge30_U0.bipedge_stream6_blk_n) | (~load_bipedge30_U0.bipedge_size_out6_blk_n);
    assign proc_1_data_PIPO_blk[7] = 1'b0;
    assign proc_1_start_FIFO_blk[7] = 1'b0;
    assign proc_1_TLF_FIFO_blk[7] = 1'b0;
    assign proc_1_input_sync_blk[7] = 1'b0 | (ap_sync_load_bipedge30_U0_ap_ready & load_bipedge30_U0.ap_idle & ~ap_sync_load_value38_U0_ap_ready);
    assign proc_1_output_sync_blk[7] = 1'b0;
    assign proc_dep_vld_vec_1[7] = dl_detect_out ? proc_dep_vld_vec_1_reg[7] : (proc_1_data_FIFO_blk[7] | proc_1_data_PIPO_blk[7] | proc_1_start_FIFO_blk[7] | proc_1_TLF_FIFO_blk[7] | proc_1_input_sync_blk[7] | proc_1_output_sync_blk[7]);
    assign proc_1_data_FIFO_blk[8] = 1'b0 | (~load_bipedge30_U0.bipedge_stream7_blk_n) | (~load_bipedge30_U0.bipedge_size_out7_blk_n);
    assign proc_1_data_PIPO_blk[8] = 1'b0;
    assign proc_1_start_FIFO_blk[8] = 1'b0;
    assign proc_1_TLF_FIFO_blk[8] = 1'b0;
    assign proc_1_input_sync_blk[8] = 1'b0 | (ap_sync_load_bipedge30_U0_ap_ready & load_bipedge30_U0.ap_idle & ~ap_sync_load_value39_U0_ap_ready);
    assign proc_1_output_sync_blk[8] = 1'b0;
    assign proc_dep_vld_vec_1[8] = dl_detect_out ? proc_dep_vld_vec_1_reg[8] : (proc_1_data_FIFO_blk[8] | proc_1_data_PIPO_blk[8] | proc_1_start_FIFO_blk[8] | proc_1_TLF_FIFO_blk[8] | proc_1_input_sync_blk[8] | proc_1_output_sync_blk[8]);
    assign proc_1_data_FIFO_blk[9] = 1'b0;
    assign proc_1_data_PIPO_blk[9] = 1'b0;
    assign proc_1_start_FIFO_blk[9] = 1'b0;
    assign proc_1_TLF_FIFO_blk[9] = 1'b0;
    assign proc_1_input_sync_blk[9] = 1'b0 | (ap_sync_load_bipedge30_U0_ap_ready & load_bipedge30_U0.ap_idle & ~ap_sync_load_bipedge31_U0_ap_ready);
    assign proc_1_output_sync_blk[9] = 1'b0;
    assign proc_dep_vld_vec_1[9] = dl_detect_out ? proc_dep_vld_vec_1_reg[9] : (proc_1_data_FIFO_blk[9] | proc_1_data_PIPO_blk[9] | proc_1_start_FIFO_blk[9] | proc_1_TLF_FIFO_blk[9] | proc_1_input_sync_blk[9] | proc_1_output_sync_blk[9]);
    assign proc_1_data_FIFO_blk[10] = 1'b0;
    assign proc_1_data_PIPO_blk[10] = 1'b0;
    assign proc_1_start_FIFO_blk[10] = 1'b0;
    assign proc_1_TLF_FIFO_blk[10] = 1'b0;
    assign proc_1_input_sync_blk[10] = 1'b0 | (ap_sync_load_bipedge30_U0_ap_ready & load_bipedge30_U0.ap_idle & ~ap_sync_load_value40_U0_ap_ready);
    assign proc_1_output_sync_blk[10] = 1'b0;
    assign proc_dep_vld_vec_1[10] = dl_detect_out ? proc_dep_vld_vec_1_reg[10] : (proc_1_data_FIFO_blk[10] | proc_1_data_PIPO_blk[10] | proc_1_start_FIFO_blk[10] | proc_1_TLF_FIFO_blk[10] | proc_1_input_sync_blk[10] | proc_1_output_sync_blk[10]);
    assign proc_1_data_FIFO_blk[11] = 1'b0;
    assign proc_1_data_PIPO_blk[11] = 1'b0;
    assign proc_1_start_FIFO_blk[11] = 1'b0;
    assign proc_1_TLF_FIFO_blk[11] = 1'b0;
    assign proc_1_input_sync_blk[11] = 1'b0 | (ap_sync_load_bipedge30_U0_ap_ready & load_bipedge30_U0.ap_idle & ~ap_sync_load_value41_U0_ap_ready);
    assign proc_1_output_sync_blk[11] = 1'b0;
    assign proc_dep_vld_vec_1[11] = dl_detect_out ? proc_dep_vld_vec_1_reg[11] : (proc_1_data_FIFO_blk[11] | proc_1_data_PIPO_blk[11] | proc_1_start_FIFO_blk[11] | proc_1_TLF_FIFO_blk[11] | proc_1_input_sync_blk[11] | proc_1_output_sync_blk[11]);
    assign proc_1_data_FIFO_blk[12] = 1'b0;
    assign proc_1_data_PIPO_blk[12] = 1'b0;
    assign proc_1_start_FIFO_blk[12] = 1'b0;
    assign proc_1_TLF_FIFO_blk[12] = 1'b0;
    assign proc_1_input_sync_blk[12] = 1'b0 | (ap_sync_load_bipedge30_U0_ap_ready & load_bipedge30_U0.ap_idle & ~ap_sync_load_value42_U0_ap_ready);
    assign proc_1_output_sync_blk[12] = 1'b0;
    assign proc_dep_vld_vec_1[12] = dl_detect_out ? proc_dep_vld_vec_1_reg[12] : (proc_1_data_FIFO_blk[12] | proc_1_data_PIPO_blk[12] | proc_1_start_FIFO_blk[12] | proc_1_TLF_FIFO_blk[12] | proc_1_input_sync_blk[12] | proc_1_output_sync_blk[12]);
    assign proc_1_data_FIFO_blk[13] = 1'b0;
    assign proc_1_data_PIPO_blk[13] = 1'b0;
    assign proc_1_start_FIFO_blk[13] = 1'b0;
    assign proc_1_TLF_FIFO_blk[13] = 1'b0;
    assign proc_1_input_sync_blk[13] = 1'b0 | (ap_sync_load_bipedge30_U0_ap_ready & load_bipedge30_U0.ap_idle & ~ap_sync_load_value43_U0_ap_ready);
    assign proc_1_output_sync_blk[13] = 1'b0;
    assign proc_dep_vld_vec_1[13] = dl_detect_out ? proc_dep_vld_vec_1_reg[13] : (proc_1_data_FIFO_blk[13] | proc_1_data_PIPO_blk[13] | proc_1_start_FIFO_blk[13] | proc_1_TLF_FIFO_blk[13] | proc_1_input_sync_blk[13] | proc_1_output_sync_blk[13]);
    assign proc_1_data_FIFO_blk[14] = 1'b0;
    assign proc_1_data_PIPO_blk[14] = 1'b0;
    assign proc_1_start_FIFO_blk[14] = 1'b0;
    assign proc_1_TLF_FIFO_blk[14] = 1'b0;
    assign proc_1_input_sync_blk[14] = 1'b0 | (ap_sync_load_bipedge30_U0_ap_ready & load_bipedge30_U0.ap_idle & ~ap_sync_load_value44_U0_ap_ready);
    assign proc_1_output_sync_blk[14] = 1'b0;
    assign proc_dep_vld_vec_1[14] = dl_detect_out ? proc_dep_vld_vec_1_reg[14] : (proc_1_data_FIFO_blk[14] | proc_1_data_PIPO_blk[14] | proc_1_start_FIFO_blk[14] | proc_1_TLF_FIFO_blk[14] | proc_1_input_sync_blk[14] | proc_1_output_sync_blk[14]);
    assign proc_1_data_FIFO_blk[15] = 1'b0;
    assign proc_1_data_PIPO_blk[15] = 1'b0;
    assign proc_1_start_FIFO_blk[15] = 1'b0;
    assign proc_1_TLF_FIFO_blk[15] = 1'b0;
    assign proc_1_input_sync_blk[15] = 1'b0 | (ap_sync_load_bipedge30_U0_ap_ready & load_bipedge30_U0.ap_idle & ~ap_sync_load_value45_U0_ap_ready);
    assign proc_1_output_sync_blk[15] = 1'b0;
    assign proc_dep_vld_vec_1[15] = dl_detect_out ? proc_dep_vld_vec_1_reg[15] : (proc_1_data_FIFO_blk[15] | proc_1_data_PIPO_blk[15] | proc_1_start_FIFO_blk[15] | proc_1_TLF_FIFO_blk[15] | proc_1_input_sync_blk[15] | proc_1_output_sync_blk[15]);
    assign proc_1_data_FIFO_blk[16] = 1'b0;
    assign proc_1_data_PIPO_blk[16] = 1'b0;
    assign proc_1_start_FIFO_blk[16] = 1'b0;
    assign proc_1_TLF_FIFO_blk[16] = 1'b0;
    assign proc_1_input_sync_blk[16] = 1'b0 | (ap_sync_load_bipedge30_U0_ap_ready & load_bipedge30_U0.ap_idle & ~ap_sync_load_value46_U0_ap_ready);
    assign proc_1_output_sync_blk[16] = 1'b0;
    assign proc_dep_vld_vec_1[16] = dl_detect_out ? proc_dep_vld_vec_1_reg[16] : (proc_1_data_FIFO_blk[16] | proc_1_data_PIPO_blk[16] | proc_1_start_FIFO_blk[16] | proc_1_TLF_FIFO_blk[16] | proc_1_input_sync_blk[16] | proc_1_output_sync_blk[16]);
    assign proc_1_data_FIFO_blk[17] = 1'b0;
    assign proc_1_data_PIPO_blk[17] = 1'b0;
    assign proc_1_start_FIFO_blk[17] = 1'b0;
    assign proc_1_TLF_FIFO_blk[17] = 1'b0;
    assign proc_1_input_sync_blk[17] = 1'b0 | (ap_sync_load_bipedge30_U0_ap_ready & load_bipedge30_U0.ap_idle & ~ap_sync_load_value47_U0_ap_ready);
    assign proc_1_output_sync_blk[17] = 1'b0;
    assign proc_dep_vld_vec_1[17] = dl_detect_out ? proc_dep_vld_vec_1_reg[17] : (proc_1_data_FIFO_blk[17] | proc_1_data_PIPO_blk[17] | proc_1_start_FIFO_blk[17] | proc_1_TLF_FIFO_blk[17] | proc_1_input_sync_blk[17] | proc_1_output_sync_blk[17]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_1_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_1_reg <= proc_dep_vld_vec_1;
        end
    end
    assign in_chan_dep_vld_vec_1[0] = dep_chan_vld_0_1;
    assign in_chan_dep_data_vec_1[34 : 0] = dep_chan_data_0_1;
    assign token_in_vec_1[0] = token_0_1;
    assign in_chan_dep_vld_vec_1[1] = dep_chan_vld_2_1;
    assign in_chan_dep_data_vec_1[69 : 35] = dep_chan_data_2_1;
    assign token_in_vec_1[1] = token_2_1;
    assign in_chan_dep_vld_vec_1[2] = dep_chan_vld_3_1;
    assign in_chan_dep_data_vec_1[104 : 70] = dep_chan_data_3_1;
    assign token_in_vec_1[2] = token_3_1;
    assign in_chan_dep_vld_vec_1[3] = dep_chan_vld_4_1;
    assign in_chan_dep_data_vec_1[139 : 105] = dep_chan_data_4_1;
    assign token_in_vec_1[3] = token_4_1;
    assign in_chan_dep_vld_vec_1[4] = dep_chan_vld_5_1;
    assign in_chan_dep_data_vec_1[174 : 140] = dep_chan_data_5_1;
    assign token_in_vec_1[4] = token_5_1;
    assign in_chan_dep_vld_vec_1[5] = dep_chan_vld_6_1;
    assign in_chan_dep_data_vec_1[209 : 175] = dep_chan_data_6_1;
    assign token_in_vec_1[5] = token_6_1;
    assign in_chan_dep_vld_vec_1[6] = dep_chan_vld_7_1;
    assign in_chan_dep_data_vec_1[244 : 210] = dep_chan_data_7_1;
    assign token_in_vec_1[6] = token_7_1;
    assign in_chan_dep_vld_vec_1[7] = dep_chan_vld_8_1;
    assign in_chan_dep_data_vec_1[279 : 245] = dep_chan_data_8_1;
    assign token_in_vec_1[7] = token_8_1;
    assign in_chan_dep_vld_vec_1[8] = dep_chan_vld_9_1;
    assign in_chan_dep_data_vec_1[314 : 280] = dep_chan_data_9_1;
    assign token_in_vec_1[8] = token_9_1;
    assign in_chan_dep_vld_vec_1[9] = dep_chan_vld_10_1;
    assign in_chan_dep_data_vec_1[349 : 315] = dep_chan_data_10_1;
    assign token_in_vec_1[9] = token_10_1;
    assign in_chan_dep_vld_vec_1[10] = dep_chan_vld_11_1;
    assign in_chan_dep_data_vec_1[384 : 350] = dep_chan_data_11_1;
    assign token_in_vec_1[10] = token_11_1;
    assign in_chan_dep_vld_vec_1[11] = dep_chan_vld_12_1;
    assign in_chan_dep_data_vec_1[419 : 385] = dep_chan_data_12_1;
    assign token_in_vec_1[11] = token_12_1;
    assign in_chan_dep_vld_vec_1[12] = dep_chan_vld_13_1;
    assign in_chan_dep_data_vec_1[454 : 420] = dep_chan_data_13_1;
    assign token_in_vec_1[12] = token_13_1;
    assign in_chan_dep_vld_vec_1[13] = dep_chan_vld_14_1;
    assign in_chan_dep_data_vec_1[489 : 455] = dep_chan_data_14_1;
    assign token_in_vec_1[13] = token_14_1;
    assign in_chan_dep_vld_vec_1[14] = dep_chan_vld_15_1;
    assign in_chan_dep_data_vec_1[524 : 490] = dep_chan_data_15_1;
    assign token_in_vec_1[14] = token_15_1;
    assign in_chan_dep_vld_vec_1[15] = dep_chan_vld_16_1;
    assign in_chan_dep_data_vec_1[559 : 525] = dep_chan_data_16_1;
    assign token_in_vec_1[15] = token_16_1;
    assign in_chan_dep_vld_vec_1[16] = dep_chan_vld_17_1;
    assign in_chan_dep_data_vec_1[594 : 560] = dep_chan_data_17_1;
    assign token_in_vec_1[16] = token_17_1;
    assign in_chan_dep_vld_vec_1[17] = dep_chan_vld_18_1;
    assign in_chan_dep_data_vec_1[629 : 595] = dep_chan_data_18_1;
    assign token_in_vec_1[17] = token_18_1;
    assign dep_chan_vld_1_0 = out_chan_dep_vld_vec_1[0];
    assign dep_chan_data_1_0 = out_chan_dep_data_1;
    assign token_1_0 = token_out_vec_1[0];
    assign dep_chan_vld_1_3 = out_chan_dep_vld_vec_1[1];
    assign dep_chan_data_1_3 = out_chan_dep_data_1;
    assign token_1_3 = token_out_vec_1[1];
    assign dep_chan_vld_1_4 = out_chan_dep_vld_vec_1[2];
    assign dep_chan_data_1_4 = out_chan_dep_data_1;
    assign token_1_4 = token_out_vec_1[2];
    assign dep_chan_vld_1_5 = out_chan_dep_vld_vec_1[3];
    assign dep_chan_data_1_5 = out_chan_dep_data_1;
    assign token_1_5 = token_out_vec_1[3];
    assign dep_chan_vld_1_6 = out_chan_dep_vld_vec_1[4];
    assign dep_chan_data_1_6 = out_chan_dep_data_1;
    assign token_1_6 = token_out_vec_1[4];
    assign dep_chan_vld_1_7 = out_chan_dep_vld_vec_1[5];
    assign dep_chan_data_1_7 = out_chan_dep_data_1;
    assign token_1_7 = token_out_vec_1[5];
    assign dep_chan_vld_1_8 = out_chan_dep_vld_vec_1[6];
    assign dep_chan_data_1_8 = out_chan_dep_data_1;
    assign token_1_8 = token_out_vec_1[6];
    assign dep_chan_vld_1_9 = out_chan_dep_vld_vec_1[7];
    assign dep_chan_data_1_9 = out_chan_dep_data_1;
    assign token_1_9 = token_out_vec_1[7];
    assign dep_chan_vld_1_10 = out_chan_dep_vld_vec_1[8];
    assign dep_chan_data_1_10 = out_chan_dep_data_1;
    assign token_1_10 = token_out_vec_1[8];
    assign dep_chan_vld_1_2 = out_chan_dep_vld_vec_1[9];
    assign dep_chan_data_1_2 = out_chan_dep_data_1;
    assign token_1_2 = token_out_vec_1[9];
    assign dep_chan_vld_1_11 = out_chan_dep_vld_vec_1[10];
    assign dep_chan_data_1_11 = out_chan_dep_data_1;
    assign token_1_11 = token_out_vec_1[10];
    assign dep_chan_vld_1_12 = out_chan_dep_vld_vec_1[11];
    assign dep_chan_data_1_12 = out_chan_dep_data_1;
    assign token_1_12 = token_out_vec_1[11];
    assign dep_chan_vld_1_13 = out_chan_dep_vld_vec_1[12];
    assign dep_chan_data_1_13 = out_chan_dep_data_1;
    assign token_1_13 = token_out_vec_1[12];
    assign dep_chan_vld_1_14 = out_chan_dep_vld_vec_1[13];
    assign dep_chan_data_1_14 = out_chan_dep_data_1;
    assign token_1_14 = token_out_vec_1[13];
    assign dep_chan_vld_1_15 = out_chan_dep_vld_vec_1[14];
    assign dep_chan_data_1_15 = out_chan_dep_data_1;
    assign token_1_15 = token_out_vec_1[14];
    assign dep_chan_vld_1_16 = out_chan_dep_vld_vec_1[15];
    assign dep_chan_data_1_16 = out_chan_dep_data_1;
    assign token_1_16 = token_out_vec_1[15];
    assign dep_chan_vld_1_17 = out_chan_dep_vld_vec_1[16];
    assign dep_chan_data_1_17 = out_chan_dep_data_1;
    assign token_1_17 = token_out_vec_1[16];
    assign dep_chan_vld_1_18 = out_chan_dep_vld_vec_1[17];
    assign dep_chan_data_1_18 = out_chan_dep_data_1;
    assign token_1_18 = token_out_vec_1[17];

    // Process: load_bipedge31_U0
    kernel_pr_hls_deadlock_detect_unit #(35, 2, 18, 18) kernel_pr_hls_deadlock_detect_unit_2 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_2),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_2),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_2),
        .token_in_vec(token_in_vec_2),
        .dl_detect_in(dl_detect_out),
        .origin(origin[2]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_2),
        .out_chan_dep_data(out_chan_dep_data_2),
        .token_out_vec(token_out_vec_2),
        .dl_detect_out(dl_in_vec[2]));

    assign proc_2_data_FIFO_blk[0] = 1'b0 | (~load_bipedge31_U0.bipedge_blk_n) | (~load_bipedge31_U0.bipedge_size_blk_n);
    assign proc_2_data_PIPO_blk[0] = 1'b0;
    assign proc_2_start_FIFO_blk[0] = 1'b0;
    assign proc_2_TLF_FIFO_blk[0] = 1'b0;
    assign proc_2_input_sync_blk[0] = 1'b0 | (ap_sync_load_bipedge31_U0_ap_ready & load_bipedge31_U0.ap_idle & ~ap_sync_kernel_pr_entry98_U0_ap_ready);
    assign proc_2_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_2[0] = dl_detect_out ? proc_dep_vld_vec_2_reg[0] : (proc_2_data_FIFO_blk[0] | proc_2_data_PIPO_blk[0] | proc_2_start_FIFO_blk[0] | proc_2_TLF_FIFO_blk[0] | proc_2_input_sync_blk[0] | proc_2_output_sync_blk[0]);
    assign proc_2_data_FIFO_blk[1] = 1'b0 | (~load_bipedge31_U0.bipedge_stream8_blk_n) | (~load_bipedge31_U0.bipedge_size_out_blk_n);
    assign proc_2_data_PIPO_blk[1] = 1'b0;
    assign proc_2_start_FIFO_blk[1] = 1'b0;
    assign proc_2_TLF_FIFO_blk[1] = 1'b0;
    assign proc_2_input_sync_blk[1] = 1'b0 | (ap_sync_load_bipedge31_U0_ap_ready & load_bipedge31_U0.ap_idle & ~ap_sync_load_value40_U0_ap_ready);
    assign proc_2_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_2[1] = dl_detect_out ? proc_dep_vld_vec_2_reg[1] : (proc_2_data_FIFO_blk[1] | proc_2_data_PIPO_blk[1] | proc_2_start_FIFO_blk[1] | proc_2_TLF_FIFO_blk[1] | proc_2_input_sync_blk[1] | proc_2_output_sync_blk[1]);
    assign proc_2_data_FIFO_blk[2] = 1'b0 | (~load_bipedge31_U0.bipedge_stream9_blk_n) | (~load_bipedge31_U0.bipedge_size_out1_blk_n);
    assign proc_2_data_PIPO_blk[2] = 1'b0;
    assign proc_2_start_FIFO_blk[2] = 1'b0;
    assign proc_2_TLF_FIFO_blk[2] = 1'b0;
    assign proc_2_input_sync_blk[2] = 1'b0 | (ap_sync_load_bipedge31_U0_ap_ready & load_bipedge31_U0.ap_idle & ~ap_sync_load_value41_U0_ap_ready);
    assign proc_2_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_2[2] = dl_detect_out ? proc_dep_vld_vec_2_reg[2] : (proc_2_data_FIFO_blk[2] | proc_2_data_PIPO_blk[2] | proc_2_start_FIFO_blk[2] | proc_2_TLF_FIFO_blk[2] | proc_2_input_sync_blk[2] | proc_2_output_sync_blk[2]);
    assign proc_2_data_FIFO_blk[3] = 1'b0 | (~load_bipedge31_U0.bipedge_stream10_blk_n) | (~load_bipedge31_U0.bipedge_size_out2_blk_n);
    assign proc_2_data_PIPO_blk[3] = 1'b0;
    assign proc_2_start_FIFO_blk[3] = 1'b0;
    assign proc_2_TLF_FIFO_blk[3] = 1'b0;
    assign proc_2_input_sync_blk[3] = 1'b0 | (ap_sync_load_bipedge31_U0_ap_ready & load_bipedge31_U0.ap_idle & ~ap_sync_load_value42_U0_ap_ready);
    assign proc_2_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_2[3] = dl_detect_out ? proc_dep_vld_vec_2_reg[3] : (proc_2_data_FIFO_blk[3] | proc_2_data_PIPO_blk[3] | proc_2_start_FIFO_blk[3] | proc_2_TLF_FIFO_blk[3] | proc_2_input_sync_blk[3] | proc_2_output_sync_blk[3]);
    assign proc_2_data_FIFO_blk[4] = 1'b0 | (~load_bipedge31_U0.bipedge_stream11_blk_n) | (~load_bipedge31_U0.bipedge_size_out3_blk_n);
    assign proc_2_data_PIPO_blk[4] = 1'b0;
    assign proc_2_start_FIFO_blk[4] = 1'b0;
    assign proc_2_TLF_FIFO_blk[4] = 1'b0;
    assign proc_2_input_sync_blk[4] = 1'b0 | (ap_sync_load_bipedge31_U0_ap_ready & load_bipedge31_U0.ap_idle & ~ap_sync_load_value43_U0_ap_ready);
    assign proc_2_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_2[4] = dl_detect_out ? proc_dep_vld_vec_2_reg[4] : (proc_2_data_FIFO_blk[4] | proc_2_data_PIPO_blk[4] | proc_2_start_FIFO_blk[4] | proc_2_TLF_FIFO_blk[4] | proc_2_input_sync_blk[4] | proc_2_output_sync_blk[4]);
    assign proc_2_data_FIFO_blk[5] = 1'b0 | (~load_bipedge31_U0.bipedge_stream12_blk_n) | (~load_bipedge31_U0.bipedge_size_out4_blk_n);
    assign proc_2_data_PIPO_blk[5] = 1'b0;
    assign proc_2_start_FIFO_blk[5] = 1'b0;
    assign proc_2_TLF_FIFO_blk[5] = 1'b0;
    assign proc_2_input_sync_blk[5] = 1'b0 | (ap_sync_load_bipedge31_U0_ap_ready & load_bipedge31_U0.ap_idle & ~ap_sync_load_value44_U0_ap_ready);
    assign proc_2_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_2[5] = dl_detect_out ? proc_dep_vld_vec_2_reg[5] : (proc_2_data_FIFO_blk[5] | proc_2_data_PIPO_blk[5] | proc_2_start_FIFO_blk[5] | proc_2_TLF_FIFO_blk[5] | proc_2_input_sync_blk[5] | proc_2_output_sync_blk[5]);
    assign proc_2_data_FIFO_blk[6] = 1'b0 | (~load_bipedge31_U0.bipedge_stream13_blk_n) | (~load_bipedge31_U0.bipedge_size_out5_blk_n);
    assign proc_2_data_PIPO_blk[6] = 1'b0;
    assign proc_2_start_FIFO_blk[6] = 1'b0;
    assign proc_2_TLF_FIFO_blk[6] = 1'b0;
    assign proc_2_input_sync_blk[6] = 1'b0 | (ap_sync_load_bipedge31_U0_ap_ready & load_bipedge31_U0.ap_idle & ~ap_sync_load_value45_U0_ap_ready);
    assign proc_2_output_sync_blk[6] = 1'b0;
    assign proc_dep_vld_vec_2[6] = dl_detect_out ? proc_dep_vld_vec_2_reg[6] : (proc_2_data_FIFO_blk[6] | proc_2_data_PIPO_blk[6] | proc_2_start_FIFO_blk[6] | proc_2_TLF_FIFO_blk[6] | proc_2_input_sync_blk[6] | proc_2_output_sync_blk[6]);
    assign proc_2_data_FIFO_blk[7] = 1'b0 | (~load_bipedge31_U0.bipedge_stream14_blk_n) | (~load_bipedge31_U0.bipedge_size_out6_blk_n);
    assign proc_2_data_PIPO_blk[7] = 1'b0;
    assign proc_2_start_FIFO_blk[7] = 1'b0;
    assign proc_2_TLF_FIFO_blk[7] = 1'b0;
    assign proc_2_input_sync_blk[7] = 1'b0 | (ap_sync_load_bipedge31_U0_ap_ready & load_bipedge31_U0.ap_idle & ~ap_sync_load_value46_U0_ap_ready);
    assign proc_2_output_sync_blk[7] = 1'b0;
    assign proc_dep_vld_vec_2[7] = dl_detect_out ? proc_dep_vld_vec_2_reg[7] : (proc_2_data_FIFO_blk[7] | proc_2_data_PIPO_blk[7] | proc_2_start_FIFO_blk[7] | proc_2_TLF_FIFO_blk[7] | proc_2_input_sync_blk[7] | proc_2_output_sync_blk[7]);
    assign proc_2_data_FIFO_blk[8] = 1'b0 | (~load_bipedge31_U0.bipedge_stream15_blk_n) | (~load_bipedge31_U0.bipedge_size_out7_blk_n);
    assign proc_2_data_PIPO_blk[8] = 1'b0;
    assign proc_2_start_FIFO_blk[8] = 1'b0;
    assign proc_2_TLF_FIFO_blk[8] = 1'b0;
    assign proc_2_input_sync_blk[8] = 1'b0 | (ap_sync_load_bipedge31_U0_ap_ready & load_bipedge31_U0.ap_idle & ~ap_sync_load_value47_U0_ap_ready);
    assign proc_2_output_sync_blk[8] = 1'b0;
    assign proc_dep_vld_vec_2[8] = dl_detect_out ? proc_dep_vld_vec_2_reg[8] : (proc_2_data_FIFO_blk[8] | proc_2_data_PIPO_blk[8] | proc_2_start_FIFO_blk[8] | proc_2_TLF_FIFO_blk[8] | proc_2_input_sync_blk[8] | proc_2_output_sync_blk[8]);
    assign proc_2_data_FIFO_blk[9] = 1'b0;
    assign proc_2_data_PIPO_blk[9] = 1'b0;
    assign proc_2_start_FIFO_blk[9] = 1'b0;
    assign proc_2_TLF_FIFO_blk[9] = 1'b0;
    assign proc_2_input_sync_blk[9] = 1'b0 | (ap_sync_load_bipedge31_U0_ap_ready & load_bipedge31_U0.ap_idle & ~ap_sync_load_bipedge30_U0_ap_ready);
    assign proc_2_output_sync_blk[9] = 1'b0;
    assign proc_dep_vld_vec_2[9] = dl_detect_out ? proc_dep_vld_vec_2_reg[9] : (proc_2_data_FIFO_blk[9] | proc_2_data_PIPO_blk[9] | proc_2_start_FIFO_blk[9] | proc_2_TLF_FIFO_blk[9] | proc_2_input_sync_blk[9] | proc_2_output_sync_blk[9]);
    assign proc_2_data_FIFO_blk[10] = 1'b0;
    assign proc_2_data_PIPO_blk[10] = 1'b0;
    assign proc_2_start_FIFO_blk[10] = 1'b0;
    assign proc_2_TLF_FIFO_blk[10] = 1'b0;
    assign proc_2_input_sync_blk[10] = 1'b0 | (ap_sync_load_bipedge31_U0_ap_ready & load_bipedge31_U0.ap_idle & ~ap_sync_load_value32_U0_ap_ready);
    assign proc_2_output_sync_blk[10] = 1'b0;
    assign proc_dep_vld_vec_2[10] = dl_detect_out ? proc_dep_vld_vec_2_reg[10] : (proc_2_data_FIFO_blk[10] | proc_2_data_PIPO_blk[10] | proc_2_start_FIFO_blk[10] | proc_2_TLF_FIFO_blk[10] | proc_2_input_sync_blk[10] | proc_2_output_sync_blk[10]);
    assign proc_2_data_FIFO_blk[11] = 1'b0;
    assign proc_2_data_PIPO_blk[11] = 1'b0;
    assign proc_2_start_FIFO_blk[11] = 1'b0;
    assign proc_2_TLF_FIFO_blk[11] = 1'b0;
    assign proc_2_input_sync_blk[11] = 1'b0 | (ap_sync_load_bipedge31_U0_ap_ready & load_bipedge31_U0.ap_idle & ~ap_sync_load_value33_U0_ap_ready);
    assign proc_2_output_sync_blk[11] = 1'b0;
    assign proc_dep_vld_vec_2[11] = dl_detect_out ? proc_dep_vld_vec_2_reg[11] : (proc_2_data_FIFO_blk[11] | proc_2_data_PIPO_blk[11] | proc_2_start_FIFO_blk[11] | proc_2_TLF_FIFO_blk[11] | proc_2_input_sync_blk[11] | proc_2_output_sync_blk[11]);
    assign proc_2_data_FIFO_blk[12] = 1'b0;
    assign proc_2_data_PIPO_blk[12] = 1'b0;
    assign proc_2_start_FIFO_blk[12] = 1'b0;
    assign proc_2_TLF_FIFO_blk[12] = 1'b0;
    assign proc_2_input_sync_blk[12] = 1'b0 | (ap_sync_load_bipedge31_U0_ap_ready & load_bipedge31_U0.ap_idle & ~ap_sync_load_value34_U0_ap_ready);
    assign proc_2_output_sync_blk[12] = 1'b0;
    assign proc_dep_vld_vec_2[12] = dl_detect_out ? proc_dep_vld_vec_2_reg[12] : (proc_2_data_FIFO_blk[12] | proc_2_data_PIPO_blk[12] | proc_2_start_FIFO_blk[12] | proc_2_TLF_FIFO_blk[12] | proc_2_input_sync_blk[12] | proc_2_output_sync_blk[12]);
    assign proc_2_data_FIFO_blk[13] = 1'b0;
    assign proc_2_data_PIPO_blk[13] = 1'b0;
    assign proc_2_start_FIFO_blk[13] = 1'b0;
    assign proc_2_TLF_FIFO_blk[13] = 1'b0;
    assign proc_2_input_sync_blk[13] = 1'b0 | (ap_sync_load_bipedge31_U0_ap_ready & load_bipedge31_U0.ap_idle & ~ap_sync_load_value35_U0_ap_ready);
    assign proc_2_output_sync_blk[13] = 1'b0;
    assign proc_dep_vld_vec_2[13] = dl_detect_out ? proc_dep_vld_vec_2_reg[13] : (proc_2_data_FIFO_blk[13] | proc_2_data_PIPO_blk[13] | proc_2_start_FIFO_blk[13] | proc_2_TLF_FIFO_blk[13] | proc_2_input_sync_blk[13] | proc_2_output_sync_blk[13]);
    assign proc_2_data_FIFO_blk[14] = 1'b0;
    assign proc_2_data_PIPO_blk[14] = 1'b0;
    assign proc_2_start_FIFO_blk[14] = 1'b0;
    assign proc_2_TLF_FIFO_blk[14] = 1'b0;
    assign proc_2_input_sync_blk[14] = 1'b0 | (ap_sync_load_bipedge31_U0_ap_ready & load_bipedge31_U0.ap_idle & ~ap_sync_load_value36_U0_ap_ready);
    assign proc_2_output_sync_blk[14] = 1'b0;
    assign proc_dep_vld_vec_2[14] = dl_detect_out ? proc_dep_vld_vec_2_reg[14] : (proc_2_data_FIFO_blk[14] | proc_2_data_PIPO_blk[14] | proc_2_start_FIFO_blk[14] | proc_2_TLF_FIFO_blk[14] | proc_2_input_sync_blk[14] | proc_2_output_sync_blk[14]);
    assign proc_2_data_FIFO_blk[15] = 1'b0;
    assign proc_2_data_PIPO_blk[15] = 1'b0;
    assign proc_2_start_FIFO_blk[15] = 1'b0;
    assign proc_2_TLF_FIFO_blk[15] = 1'b0;
    assign proc_2_input_sync_blk[15] = 1'b0 | (ap_sync_load_bipedge31_U0_ap_ready & load_bipedge31_U0.ap_idle & ~ap_sync_load_value37_U0_ap_ready);
    assign proc_2_output_sync_blk[15] = 1'b0;
    assign proc_dep_vld_vec_2[15] = dl_detect_out ? proc_dep_vld_vec_2_reg[15] : (proc_2_data_FIFO_blk[15] | proc_2_data_PIPO_blk[15] | proc_2_start_FIFO_blk[15] | proc_2_TLF_FIFO_blk[15] | proc_2_input_sync_blk[15] | proc_2_output_sync_blk[15]);
    assign proc_2_data_FIFO_blk[16] = 1'b0;
    assign proc_2_data_PIPO_blk[16] = 1'b0;
    assign proc_2_start_FIFO_blk[16] = 1'b0;
    assign proc_2_TLF_FIFO_blk[16] = 1'b0;
    assign proc_2_input_sync_blk[16] = 1'b0 | (ap_sync_load_bipedge31_U0_ap_ready & load_bipedge31_U0.ap_idle & ~ap_sync_load_value38_U0_ap_ready);
    assign proc_2_output_sync_blk[16] = 1'b0;
    assign proc_dep_vld_vec_2[16] = dl_detect_out ? proc_dep_vld_vec_2_reg[16] : (proc_2_data_FIFO_blk[16] | proc_2_data_PIPO_blk[16] | proc_2_start_FIFO_blk[16] | proc_2_TLF_FIFO_blk[16] | proc_2_input_sync_blk[16] | proc_2_output_sync_blk[16]);
    assign proc_2_data_FIFO_blk[17] = 1'b0;
    assign proc_2_data_PIPO_blk[17] = 1'b0;
    assign proc_2_start_FIFO_blk[17] = 1'b0;
    assign proc_2_TLF_FIFO_blk[17] = 1'b0;
    assign proc_2_input_sync_blk[17] = 1'b0 | (ap_sync_load_bipedge31_U0_ap_ready & load_bipedge31_U0.ap_idle & ~ap_sync_load_value39_U0_ap_ready);
    assign proc_2_output_sync_blk[17] = 1'b0;
    assign proc_dep_vld_vec_2[17] = dl_detect_out ? proc_dep_vld_vec_2_reg[17] : (proc_2_data_FIFO_blk[17] | proc_2_data_PIPO_blk[17] | proc_2_start_FIFO_blk[17] | proc_2_TLF_FIFO_blk[17] | proc_2_input_sync_blk[17] | proc_2_output_sync_blk[17]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_2_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_2_reg <= proc_dep_vld_vec_2;
        end
    end
    assign in_chan_dep_vld_vec_2[0] = dep_chan_vld_0_2;
    assign in_chan_dep_data_vec_2[34 : 0] = dep_chan_data_0_2;
    assign token_in_vec_2[0] = token_0_2;
    assign in_chan_dep_vld_vec_2[1] = dep_chan_vld_1_2;
    assign in_chan_dep_data_vec_2[69 : 35] = dep_chan_data_1_2;
    assign token_in_vec_2[1] = token_1_2;
    assign in_chan_dep_vld_vec_2[2] = dep_chan_vld_3_2;
    assign in_chan_dep_data_vec_2[104 : 70] = dep_chan_data_3_2;
    assign token_in_vec_2[2] = token_3_2;
    assign in_chan_dep_vld_vec_2[3] = dep_chan_vld_4_2;
    assign in_chan_dep_data_vec_2[139 : 105] = dep_chan_data_4_2;
    assign token_in_vec_2[3] = token_4_2;
    assign in_chan_dep_vld_vec_2[4] = dep_chan_vld_5_2;
    assign in_chan_dep_data_vec_2[174 : 140] = dep_chan_data_5_2;
    assign token_in_vec_2[4] = token_5_2;
    assign in_chan_dep_vld_vec_2[5] = dep_chan_vld_6_2;
    assign in_chan_dep_data_vec_2[209 : 175] = dep_chan_data_6_2;
    assign token_in_vec_2[5] = token_6_2;
    assign in_chan_dep_vld_vec_2[6] = dep_chan_vld_7_2;
    assign in_chan_dep_data_vec_2[244 : 210] = dep_chan_data_7_2;
    assign token_in_vec_2[6] = token_7_2;
    assign in_chan_dep_vld_vec_2[7] = dep_chan_vld_8_2;
    assign in_chan_dep_data_vec_2[279 : 245] = dep_chan_data_8_2;
    assign token_in_vec_2[7] = token_8_2;
    assign in_chan_dep_vld_vec_2[8] = dep_chan_vld_9_2;
    assign in_chan_dep_data_vec_2[314 : 280] = dep_chan_data_9_2;
    assign token_in_vec_2[8] = token_9_2;
    assign in_chan_dep_vld_vec_2[9] = dep_chan_vld_10_2;
    assign in_chan_dep_data_vec_2[349 : 315] = dep_chan_data_10_2;
    assign token_in_vec_2[9] = token_10_2;
    assign in_chan_dep_vld_vec_2[10] = dep_chan_vld_11_2;
    assign in_chan_dep_data_vec_2[384 : 350] = dep_chan_data_11_2;
    assign token_in_vec_2[10] = token_11_2;
    assign in_chan_dep_vld_vec_2[11] = dep_chan_vld_12_2;
    assign in_chan_dep_data_vec_2[419 : 385] = dep_chan_data_12_2;
    assign token_in_vec_2[11] = token_12_2;
    assign in_chan_dep_vld_vec_2[12] = dep_chan_vld_13_2;
    assign in_chan_dep_data_vec_2[454 : 420] = dep_chan_data_13_2;
    assign token_in_vec_2[12] = token_13_2;
    assign in_chan_dep_vld_vec_2[13] = dep_chan_vld_14_2;
    assign in_chan_dep_data_vec_2[489 : 455] = dep_chan_data_14_2;
    assign token_in_vec_2[13] = token_14_2;
    assign in_chan_dep_vld_vec_2[14] = dep_chan_vld_15_2;
    assign in_chan_dep_data_vec_2[524 : 490] = dep_chan_data_15_2;
    assign token_in_vec_2[14] = token_15_2;
    assign in_chan_dep_vld_vec_2[15] = dep_chan_vld_16_2;
    assign in_chan_dep_data_vec_2[559 : 525] = dep_chan_data_16_2;
    assign token_in_vec_2[15] = token_16_2;
    assign in_chan_dep_vld_vec_2[16] = dep_chan_vld_17_2;
    assign in_chan_dep_data_vec_2[594 : 560] = dep_chan_data_17_2;
    assign token_in_vec_2[16] = token_17_2;
    assign in_chan_dep_vld_vec_2[17] = dep_chan_vld_18_2;
    assign in_chan_dep_data_vec_2[629 : 595] = dep_chan_data_18_2;
    assign token_in_vec_2[17] = token_18_2;
    assign dep_chan_vld_2_0 = out_chan_dep_vld_vec_2[0];
    assign dep_chan_data_2_0 = out_chan_dep_data_2;
    assign token_2_0 = token_out_vec_2[0];
    assign dep_chan_vld_2_11 = out_chan_dep_vld_vec_2[1];
    assign dep_chan_data_2_11 = out_chan_dep_data_2;
    assign token_2_11 = token_out_vec_2[1];
    assign dep_chan_vld_2_12 = out_chan_dep_vld_vec_2[2];
    assign dep_chan_data_2_12 = out_chan_dep_data_2;
    assign token_2_12 = token_out_vec_2[2];
    assign dep_chan_vld_2_13 = out_chan_dep_vld_vec_2[3];
    assign dep_chan_data_2_13 = out_chan_dep_data_2;
    assign token_2_13 = token_out_vec_2[3];
    assign dep_chan_vld_2_14 = out_chan_dep_vld_vec_2[4];
    assign dep_chan_data_2_14 = out_chan_dep_data_2;
    assign token_2_14 = token_out_vec_2[4];
    assign dep_chan_vld_2_15 = out_chan_dep_vld_vec_2[5];
    assign dep_chan_data_2_15 = out_chan_dep_data_2;
    assign token_2_15 = token_out_vec_2[5];
    assign dep_chan_vld_2_16 = out_chan_dep_vld_vec_2[6];
    assign dep_chan_data_2_16 = out_chan_dep_data_2;
    assign token_2_16 = token_out_vec_2[6];
    assign dep_chan_vld_2_17 = out_chan_dep_vld_vec_2[7];
    assign dep_chan_data_2_17 = out_chan_dep_data_2;
    assign token_2_17 = token_out_vec_2[7];
    assign dep_chan_vld_2_18 = out_chan_dep_vld_vec_2[8];
    assign dep_chan_data_2_18 = out_chan_dep_data_2;
    assign token_2_18 = token_out_vec_2[8];
    assign dep_chan_vld_2_1 = out_chan_dep_vld_vec_2[9];
    assign dep_chan_data_2_1 = out_chan_dep_data_2;
    assign token_2_1 = token_out_vec_2[9];
    assign dep_chan_vld_2_3 = out_chan_dep_vld_vec_2[10];
    assign dep_chan_data_2_3 = out_chan_dep_data_2;
    assign token_2_3 = token_out_vec_2[10];
    assign dep_chan_vld_2_4 = out_chan_dep_vld_vec_2[11];
    assign dep_chan_data_2_4 = out_chan_dep_data_2;
    assign token_2_4 = token_out_vec_2[11];
    assign dep_chan_vld_2_5 = out_chan_dep_vld_vec_2[12];
    assign dep_chan_data_2_5 = out_chan_dep_data_2;
    assign token_2_5 = token_out_vec_2[12];
    assign dep_chan_vld_2_6 = out_chan_dep_vld_vec_2[13];
    assign dep_chan_data_2_6 = out_chan_dep_data_2;
    assign token_2_6 = token_out_vec_2[13];
    assign dep_chan_vld_2_7 = out_chan_dep_vld_vec_2[14];
    assign dep_chan_data_2_7 = out_chan_dep_data_2;
    assign token_2_7 = token_out_vec_2[14];
    assign dep_chan_vld_2_8 = out_chan_dep_vld_vec_2[15];
    assign dep_chan_data_2_8 = out_chan_dep_data_2;
    assign token_2_8 = token_out_vec_2[15];
    assign dep_chan_vld_2_9 = out_chan_dep_vld_vec_2[16];
    assign dep_chan_data_2_9 = out_chan_dep_data_2;
    assign token_2_9 = token_out_vec_2[16];
    assign dep_chan_vld_2_10 = out_chan_dep_vld_vec_2[17];
    assign dep_chan_data_2_10 = out_chan_dep_data_2;
    assign token_2_10 = token_out_vec_2[17];

    // Process: load_value32_U0
    kernel_pr_hls_deadlock_detect_unit #(35, 3, 19, 19) kernel_pr_hls_deadlock_detect_unit_3 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_3),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_3),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_3),
        .token_in_vec(token_in_vec_3),
        .dl_detect_in(dl_detect_out),
        .origin(origin[3]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_3),
        .out_chan_dep_data(out_chan_dep_data_3),
        .token_out_vec(token_out_vec_3),
        .dl_detect_out(dl_in_vec[3]));

    assign proc_3_data_FIFO_blk[0] = 1'b0 | (~load_value32_U0.value_r_blk_n);
    assign proc_3_data_PIPO_blk[0] = 1'b0;
    assign proc_3_start_FIFO_blk[0] = 1'b0;
    assign proc_3_TLF_FIFO_blk[0] = 1'b0;
    assign proc_3_input_sync_blk[0] = 1'b0 | (ap_sync_load_value32_U0_ap_ready & load_value32_U0.ap_idle & ~ap_sync_kernel_pr_entry98_U0_ap_ready);
    assign proc_3_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_3[0] = dl_detect_out ? proc_dep_vld_vec_3_reg[0] : (proc_3_data_FIFO_blk[0] | proc_3_data_PIPO_blk[0] | proc_3_start_FIFO_blk[0] | proc_3_TLF_FIFO_blk[0] | proc_3_input_sync_blk[0] | proc_3_output_sync_blk[0]);
    assign proc_3_data_FIFO_blk[1] = 1'b0 | (~load_value32_U0.bipedge_size_blk_n) | (~load_value32_U0.bipedge_stream_V_V_blk_n);
    assign proc_3_data_PIPO_blk[1] = 1'b0;
    assign proc_3_start_FIFO_blk[1] = 1'b0;
    assign proc_3_TLF_FIFO_blk[1] = 1'b0;
    assign proc_3_input_sync_blk[1] = 1'b0 | (ap_sync_load_value32_U0_ap_ready & load_value32_U0.ap_idle & ~ap_sync_load_bipedge30_U0_ap_ready);
    assign proc_3_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_3[1] = dl_detect_out ? proc_dep_vld_vec_3_reg[1] : (proc_3_data_FIFO_blk[1] | proc_3_data_PIPO_blk[1] | proc_3_start_FIFO_blk[1] | proc_3_TLF_FIFO_blk[1] | proc_3_input_sync_blk[1] | proc_3_output_sync_blk[1]);
    assign proc_3_data_FIFO_blk[2] = 1'b0 | (~load_value32_U0.value_stream_V_V_blk_n);
    assign proc_3_data_PIPO_blk[2] = 1'b0;
    assign proc_3_start_FIFO_blk[2] = 1'b0;
    assign proc_3_TLF_FIFO_blk[2] = 1'b0;
    assign proc_3_input_sync_blk[2] = 1'b0;
    assign proc_3_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_3[2] = dl_detect_out ? proc_dep_vld_vec_3_reg[2] : (proc_3_data_FIFO_blk[2] | proc_3_data_PIPO_blk[2] | proc_3_start_FIFO_blk[2] | proc_3_TLF_FIFO_blk[2] | proc_3_input_sync_blk[2] | proc_3_output_sync_blk[2]);
    assign proc_3_data_FIFO_blk[3] = 1'b0;
    assign proc_3_data_PIPO_blk[3] = 1'b0;
    assign proc_3_start_FIFO_blk[3] = 1'b0;
    assign proc_3_TLF_FIFO_blk[3] = 1'b0;
    assign proc_3_input_sync_blk[3] = 1'b0 | (ap_sync_load_value32_U0_ap_ready & load_value32_U0.ap_idle & ~ap_sync_load_bipedge31_U0_ap_ready);
    assign proc_3_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_3[3] = dl_detect_out ? proc_dep_vld_vec_3_reg[3] : (proc_3_data_FIFO_blk[3] | proc_3_data_PIPO_blk[3] | proc_3_start_FIFO_blk[3] | proc_3_TLF_FIFO_blk[3] | proc_3_input_sync_blk[3] | proc_3_output_sync_blk[3]);
    assign proc_3_data_FIFO_blk[4] = 1'b0;
    assign proc_3_data_PIPO_blk[4] = 1'b0;
    assign proc_3_start_FIFO_blk[4] = 1'b0;
    assign proc_3_TLF_FIFO_blk[4] = 1'b0;
    assign proc_3_input_sync_blk[4] = 1'b0 | (ap_sync_load_value32_U0_ap_ready & load_value32_U0.ap_idle & ~ap_sync_load_value33_U0_ap_ready);
    assign proc_3_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_3[4] = dl_detect_out ? proc_dep_vld_vec_3_reg[4] : (proc_3_data_FIFO_blk[4] | proc_3_data_PIPO_blk[4] | proc_3_start_FIFO_blk[4] | proc_3_TLF_FIFO_blk[4] | proc_3_input_sync_blk[4] | proc_3_output_sync_blk[4]);
    assign proc_3_data_FIFO_blk[5] = 1'b0;
    assign proc_3_data_PIPO_blk[5] = 1'b0;
    assign proc_3_start_FIFO_blk[5] = 1'b0;
    assign proc_3_TLF_FIFO_blk[5] = 1'b0;
    assign proc_3_input_sync_blk[5] = 1'b0 | (ap_sync_load_value32_U0_ap_ready & load_value32_U0.ap_idle & ~ap_sync_load_value34_U0_ap_ready);
    assign proc_3_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_3[5] = dl_detect_out ? proc_dep_vld_vec_3_reg[5] : (proc_3_data_FIFO_blk[5] | proc_3_data_PIPO_blk[5] | proc_3_start_FIFO_blk[5] | proc_3_TLF_FIFO_blk[5] | proc_3_input_sync_blk[5] | proc_3_output_sync_blk[5]);
    assign proc_3_data_FIFO_blk[6] = 1'b0;
    assign proc_3_data_PIPO_blk[6] = 1'b0;
    assign proc_3_start_FIFO_blk[6] = 1'b0;
    assign proc_3_TLF_FIFO_blk[6] = 1'b0;
    assign proc_3_input_sync_blk[6] = 1'b0 | (ap_sync_load_value32_U0_ap_ready & load_value32_U0.ap_idle & ~ap_sync_load_value35_U0_ap_ready);
    assign proc_3_output_sync_blk[6] = 1'b0;
    assign proc_dep_vld_vec_3[6] = dl_detect_out ? proc_dep_vld_vec_3_reg[6] : (proc_3_data_FIFO_blk[6] | proc_3_data_PIPO_blk[6] | proc_3_start_FIFO_blk[6] | proc_3_TLF_FIFO_blk[6] | proc_3_input_sync_blk[6] | proc_3_output_sync_blk[6]);
    assign proc_3_data_FIFO_blk[7] = 1'b0;
    assign proc_3_data_PIPO_blk[7] = 1'b0;
    assign proc_3_start_FIFO_blk[7] = 1'b0;
    assign proc_3_TLF_FIFO_blk[7] = 1'b0;
    assign proc_3_input_sync_blk[7] = 1'b0 | (ap_sync_load_value32_U0_ap_ready & load_value32_U0.ap_idle & ~ap_sync_load_value36_U0_ap_ready);
    assign proc_3_output_sync_blk[7] = 1'b0;
    assign proc_dep_vld_vec_3[7] = dl_detect_out ? proc_dep_vld_vec_3_reg[7] : (proc_3_data_FIFO_blk[7] | proc_3_data_PIPO_blk[7] | proc_3_start_FIFO_blk[7] | proc_3_TLF_FIFO_blk[7] | proc_3_input_sync_blk[7] | proc_3_output_sync_blk[7]);
    assign proc_3_data_FIFO_blk[8] = 1'b0;
    assign proc_3_data_PIPO_blk[8] = 1'b0;
    assign proc_3_start_FIFO_blk[8] = 1'b0;
    assign proc_3_TLF_FIFO_blk[8] = 1'b0;
    assign proc_3_input_sync_blk[8] = 1'b0 | (ap_sync_load_value32_U0_ap_ready & load_value32_U0.ap_idle & ~ap_sync_load_value37_U0_ap_ready);
    assign proc_3_output_sync_blk[8] = 1'b0;
    assign proc_dep_vld_vec_3[8] = dl_detect_out ? proc_dep_vld_vec_3_reg[8] : (proc_3_data_FIFO_blk[8] | proc_3_data_PIPO_blk[8] | proc_3_start_FIFO_blk[8] | proc_3_TLF_FIFO_blk[8] | proc_3_input_sync_blk[8] | proc_3_output_sync_blk[8]);
    assign proc_3_data_FIFO_blk[9] = 1'b0;
    assign proc_3_data_PIPO_blk[9] = 1'b0;
    assign proc_3_start_FIFO_blk[9] = 1'b0;
    assign proc_3_TLF_FIFO_blk[9] = 1'b0;
    assign proc_3_input_sync_blk[9] = 1'b0 | (ap_sync_load_value32_U0_ap_ready & load_value32_U0.ap_idle & ~ap_sync_load_value38_U0_ap_ready);
    assign proc_3_output_sync_blk[9] = 1'b0;
    assign proc_dep_vld_vec_3[9] = dl_detect_out ? proc_dep_vld_vec_3_reg[9] : (proc_3_data_FIFO_blk[9] | proc_3_data_PIPO_blk[9] | proc_3_start_FIFO_blk[9] | proc_3_TLF_FIFO_blk[9] | proc_3_input_sync_blk[9] | proc_3_output_sync_blk[9]);
    assign proc_3_data_FIFO_blk[10] = 1'b0;
    assign proc_3_data_PIPO_blk[10] = 1'b0;
    assign proc_3_start_FIFO_blk[10] = 1'b0;
    assign proc_3_TLF_FIFO_blk[10] = 1'b0;
    assign proc_3_input_sync_blk[10] = 1'b0 | (ap_sync_load_value32_U0_ap_ready & load_value32_U0.ap_idle & ~ap_sync_load_value39_U0_ap_ready);
    assign proc_3_output_sync_blk[10] = 1'b0;
    assign proc_dep_vld_vec_3[10] = dl_detect_out ? proc_dep_vld_vec_3_reg[10] : (proc_3_data_FIFO_blk[10] | proc_3_data_PIPO_blk[10] | proc_3_start_FIFO_blk[10] | proc_3_TLF_FIFO_blk[10] | proc_3_input_sync_blk[10] | proc_3_output_sync_blk[10]);
    assign proc_3_data_FIFO_blk[11] = 1'b0;
    assign proc_3_data_PIPO_blk[11] = 1'b0;
    assign proc_3_start_FIFO_blk[11] = 1'b0;
    assign proc_3_TLF_FIFO_blk[11] = 1'b0;
    assign proc_3_input_sync_blk[11] = 1'b0 | (ap_sync_load_value32_U0_ap_ready & load_value32_U0.ap_idle & ~ap_sync_load_value40_U0_ap_ready);
    assign proc_3_output_sync_blk[11] = 1'b0;
    assign proc_dep_vld_vec_3[11] = dl_detect_out ? proc_dep_vld_vec_3_reg[11] : (proc_3_data_FIFO_blk[11] | proc_3_data_PIPO_blk[11] | proc_3_start_FIFO_blk[11] | proc_3_TLF_FIFO_blk[11] | proc_3_input_sync_blk[11] | proc_3_output_sync_blk[11]);
    assign proc_3_data_FIFO_blk[12] = 1'b0;
    assign proc_3_data_PIPO_blk[12] = 1'b0;
    assign proc_3_start_FIFO_blk[12] = 1'b0;
    assign proc_3_TLF_FIFO_blk[12] = 1'b0;
    assign proc_3_input_sync_blk[12] = 1'b0 | (ap_sync_load_value32_U0_ap_ready & load_value32_U0.ap_idle & ~ap_sync_load_value41_U0_ap_ready);
    assign proc_3_output_sync_blk[12] = 1'b0;
    assign proc_dep_vld_vec_3[12] = dl_detect_out ? proc_dep_vld_vec_3_reg[12] : (proc_3_data_FIFO_blk[12] | proc_3_data_PIPO_blk[12] | proc_3_start_FIFO_blk[12] | proc_3_TLF_FIFO_blk[12] | proc_3_input_sync_blk[12] | proc_3_output_sync_blk[12]);
    assign proc_3_data_FIFO_blk[13] = 1'b0;
    assign proc_3_data_PIPO_blk[13] = 1'b0;
    assign proc_3_start_FIFO_blk[13] = 1'b0;
    assign proc_3_TLF_FIFO_blk[13] = 1'b0;
    assign proc_3_input_sync_blk[13] = 1'b0 | (ap_sync_load_value32_U0_ap_ready & load_value32_U0.ap_idle & ~ap_sync_load_value42_U0_ap_ready);
    assign proc_3_output_sync_blk[13] = 1'b0;
    assign proc_dep_vld_vec_3[13] = dl_detect_out ? proc_dep_vld_vec_3_reg[13] : (proc_3_data_FIFO_blk[13] | proc_3_data_PIPO_blk[13] | proc_3_start_FIFO_blk[13] | proc_3_TLF_FIFO_blk[13] | proc_3_input_sync_blk[13] | proc_3_output_sync_blk[13]);
    assign proc_3_data_FIFO_blk[14] = 1'b0;
    assign proc_3_data_PIPO_blk[14] = 1'b0;
    assign proc_3_start_FIFO_blk[14] = 1'b0;
    assign proc_3_TLF_FIFO_blk[14] = 1'b0;
    assign proc_3_input_sync_blk[14] = 1'b0 | (ap_sync_load_value32_U0_ap_ready & load_value32_U0.ap_idle & ~ap_sync_load_value43_U0_ap_ready);
    assign proc_3_output_sync_blk[14] = 1'b0;
    assign proc_dep_vld_vec_3[14] = dl_detect_out ? proc_dep_vld_vec_3_reg[14] : (proc_3_data_FIFO_blk[14] | proc_3_data_PIPO_blk[14] | proc_3_start_FIFO_blk[14] | proc_3_TLF_FIFO_blk[14] | proc_3_input_sync_blk[14] | proc_3_output_sync_blk[14]);
    assign proc_3_data_FIFO_blk[15] = 1'b0;
    assign proc_3_data_PIPO_blk[15] = 1'b0;
    assign proc_3_start_FIFO_blk[15] = 1'b0;
    assign proc_3_TLF_FIFO_blk[15] = 1'b0;
    assign proc_3_input_sync_blk[15] = 1'b0 | (ap_sync_load_value32_U0_ap_ready & load_value32_U0.ap_idle & ~ap_sync_load_value44_U0_ap_ready);
    assign proc_3_output_sync_blk[15] = 1'b0;
    assign proc_dep_vld_vec_3[15] = dl_detect_out ? proc_dep_vld_vec_3_reg[15] : (proc_3_data_FIFO_blk[15] | proc_3_data_PIPO_blk[15] | proc_3_start_FIFO_blk[15] | proc_3_TLF_FIFO_blk[15] | proc_3_input_sync_blk[15] | proc_3_output_sync_blk[15]);
    assign proc_3_data_FIFO_blk[16] = 1'b0;
    assign proc_3_data_PIPO_blk[16] = 1'b0;
    assign proc_3_start_FIFO_blk[16] = 1'b0;
    assign proc_3_TLF_FIFO_blk[16] = 1'b0;
    assign proc_3_input_sync_blk[16] = 1'b0 | (ap_sync_load_value32_U0_ap_ready & load_value32_U0.ap_idle & ~ap_sync_load_value45_U0_ap_ready);
    assign proc_3_output_sync_blk[16] = 1'b0;
    assign proc_dep_vld_vec_3[16] = dl_detect_out ? proc_dep_vld_vec_3_reg[16] : (proc_3_data_FIFO_blk[16] | proc_3_data_PIPO_blk[16] | proc_3_start_FIFO_blk[16] | proc_3_TLF_FIFO_blk[16] | proc_3_input_sync_blk[16] | proc_3_output_sync_blk[16]);
    assign proc_3_data_FIFO_blk[17] = 1'b0;
    assign proc_3_data_PIPO_blk[17] = 1'b0;
    assign proc_3_start_FIFO_blk[17] = 1'b0;
    assign proc_3_TLF_FIFO_blk[17] = 1'b0;
    assign proc_3_input_sync_blk[17] = 1'b0 | (ap_sync_load_value32_U0_ap_ready & load_value32_U0.ap_idle & ~ap_sync_load_value46_U0_ap_ready);
    assign proc_3_output_sync_blk[17] = 1'b0;
    assign proc_dep_vld_vec_3[17] = dl_detect_out ? proc_dep_vld_vec_3_reg[17] : (proc_3_data_FIFO_blk[17] | proc_3_data_PIPO_blk[17] | proc_3_start_FIFO_blk[17] | proc_3_TLF_FIFO_blk[17] | proc_3_input_sync_blk[17] | proc_3_output_sync_blk[17]);
    assign proc_3_data_FIFO_blk[18] = 1'b0;
    assign proc_3_data_PIPO_blk[18] = 1'b0;
    assign proc_3_start_FIFO_blk[18] = 1'b0;
    assign proc_3_TLF_FIFO_blk[18] = 1'b0;
    assign proc_3_input_sync_blk[18] = 1'b0 | (ap_sync_load_value32_U0_ap_ready & load_value32_U0.ap_idle & ~ap_sync_load_value47_U0_ap_ready);
    assign proc_3_output_sync_blk[18] = 1'b0;
    assign proc_dep_vld_vec_3[18] = dl_detect_out ? proc_dep_vld_vec_3_reg[18] : (proc_3_data_FIFO_blk[18] | proc_3_data_PIPO_blk[18] | proc_3_start_FIFO_blk[18] | proc_3_TLF_FIFO_blk[18] | proc_3_input_sync_blk[18] | proc_3_output_sync_blk[18]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_3_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_3_reg <= proc_dep_vld_vec_3;
        end
    end
    assign in_chan_dep_vld_vec_3[0] = dep_chan_vld_0_3;
    assign in_chan_dep_data_vec_3[34 : 0] = dep_chan_data_0_3;
    assign token_in_vec_3[0] = token_0_3;
    assign in_chan_dep_vld_vec_3[1] = dep_chan_vld_1_3;
    assign in_chan_dep_data_vec_3[69 : 35] = dep_chan_data_1_3;
    assign token_in_vec_3[1] = token_1_3;
    assign in_chan_dep_vld_vec_3[2] = dep_chan_vld_2_3;
    assign in_chan_dep_data_vec_3[104 : 70] = dep_chan_data_2_3;
    assign token_in_vec_3[2] = token_2_3;
    assign in_chan_dep_vld_vec_3[3] = dep_chan_vld_4_3;
    assign in_chan_dep_data_vec_3[139 : 105] = dep_chan_data_4_3;
    assign token_in_vec_3[3] = token_4_3;
    assign in_chan_dep_vld_vec_3[4] = dep_chan_vld_5_3;
    assign in_chan_dep_data_vec_3[174 : 140] = dep_chan_data_5_3;
    assign token_in_vec_3[4] = token_5_3;
    assign in_chan_dep_vld_vec_3[5] = dep_chan_vld_6_3;
    assign in_chan_dep_data_vec_3[209 : 175] = dep_chan_data_6_3;
    assign token_in_vec_3[5] = token_6_3;
    assign in_chan_dep_vld_vec_3[6] = dep_chan_vld_7_3;
    assign in_chan_dep_data_vec_3[244 : 210] = dep_chan_data_7_3;
    assign token_in_vec_3[6] = token_7_3;
    assign in_chan_dep_vld_vec_3[7] = dep_chan_vld_8_3;
    assign in_chan_dep_data_vec_3[279 : 245] = dep_chan_data_8_3;
    assign token_in_vec_3[7] = token_8_3;
    assign in_chan_dep_vld_vec_3[8] = dep_chan_vld_9_3;
    assign in_chan_dep_data_vec_3[314 : 280] = dep_chan_data_9_3;
    assign token_in_vec_3[8] = token_9_3;
    assign in_chan_dep_vld_vec_3[9] = dep_chan_vld_10_3;
    assign in_chan_dep_data_vec_3[349 : 315] = dep_chan_data_10_3;
    assign token_in_vec_3[9] = token_10_3;
    assign in_chan_dep_vld_vec_3[10] = dep_chan_vld_11_3;
    assign in_chan_dep_data_vec_3[384 : 350] = dep_chan_data_11_3;
    assign token_in_vec_3[10] = token_11_3;
    assign in_chan_dep_vld_vec_3[11] = dep_chan_vld_12_3;
    assign in_chan_dep_data_vec_3[419 : 385] = dep_chan_data_12_3;
    assign token_in_vec_3[11] = token_12_3;
    assign in_chan_dep_vld_vec_3[12] = dep_chan_vld_13_3;
    assign in_chan_dep_data_vec_3[454 : 420] = dep_chan_data_13_3;
    assign token_in_vec_3[12] = token_13_3;
    assign in_chan_dep_vld_vec_3[13] = dep_chan_vld_14_3;
    assign in_chan_dep_data_vec_3[489 : 455] = dep_chan_data_14_3;
    assign token_in_vec_3[13] = token_14_3;
    assign in_chan_dep_vld_vec_3[14] = dep_chan_vld_15_3;
    assign in_chan_dep_data_vec_3[524 : 490] = dep_chan_data_15_3;
    assign token_in_vec_3[14] = token_15_3;
    assign in_chan_dep_vld_vec_3[15] = dep_chan_vld_16_3;
    assign in_chan_dep_data_vec_3[559 : 525] = dep_chan_data_16_3;
    assign token_in_vec_3[15] = token_16_3;
    assign in_chan_dep_vld_vec_3[16] = dep_chan_vld_17_3;
    assign in_chan_dep_data_vec_3[594 : 560] = dep_chan_data_17_3;
    assign token_in_vec_3[16] = token_17_3;
    assign in_chan_dep_vld_vec_3[17] = dep_chan_vld_18_3;
    assign in_chan_dep_data_vec_3[629 : 595] = dep_chan_data_18_3;
    assign token_in_vec_3[17] = token_18_3;
    assign in_chan_dep_vld_vec_3[18] = dep_chan_vld_19_3;
    assign in_chan_dep_data_vec_3[664 : 630] = dep_chan_data_19_3;
    assign token_in_vec_3[18] = token_19_3;
    assign dep_chan_vld_3_0 = out_chan_dep_vld_vec_3[0];
    assign dep_chan_data_3_0 = out_chan_dep_data_3;
    assign token_3_0 = token_out_vec_3[0];
    assign dep_chan_vld_3_1 = out_chan_dep_vld_vec_3[1];
    assign dep_chan_data_3_1 = out_chan_dep_data_3;
    assign token_3_1 = token_out_vec_3[1];
    assign dep_chan_vld_3_19 = out_chan_dep_vld_vec_3[2];
    assign dep_chan_data_3_19 = out_chan_dep_data_3;
    assign token_3_19 = token_out_vec_3[2];
    assign dep_chan_vld_3_2 = out_chan_dep_vld_vec_3[3];
    assign dep_chan_data_3_2 = out_chan_dep_data_3;
    assign token_3_2 = token_out_vec_3[3];
    assign dep_chan_vld_3_4 = out_chan_dep_vld_vec_3[4];
    assign dep_chan_data_3_4 = out_chan_dep_data_3;
    assign token_3_4 = token_out_vec_3[4];
    assign dep_chan_vld_3_5 = out_chan_dep_vld_vec_3[5];
    assign dep_chan_data_3_5 = out_chan_dep_data_3;
    assign token_3_5 = token_out_vec_3[5];
    assign dep_chan_vld_3_6 = out_chan_dep_vld_vec_3[6];
    assign dep_chan_data_3_6 = out_chan_dep_data_3;
    assign token_3_6 = token_out_vec_3[6];
    assign dep_chan_vld_3_7 = out_chan_dep_vld_vec_3[7];
    assign dep_chan_data_3_7 = out_chan_dep_data_3;
    assign token_3_7 = token_out_vec_3[7];
    assign dep_chan_vld_3_8 = out_chan_dep_vld_vec_3[8];
    assign dep_chan_data_3_8 = out_chan_dep_data_3;
    assign token_3_8 = token_out_vec_3[8];
    assign dep_chan_vld_3_9 = out_chan_dep_vld_vec_3[9];
    assign dep_chan_data_3_9 = out_chan_dep_data_3;
    assign token_3_9 = token_out_vec_3[9];
    assign dep_chan_vld_3_10 = out_chan_dep_vld_vec_3[10];
    assign dep_chan_data_3_10 = out_chan_dep_data_3;
    assign token_3_10 = token_out_vec_3[10];
    assign dep_chan_vld_3_11 = out_chan_dep_vld_vec_3[11];
    assign dep_chan_data_3_11 = out_chan_dep_data_3;
    assign token_3_11 = token_out_vec_3[11];
    assign dep_chan_vld_3_12 = out_chan_dep_vld_vec_3[12];
    assign dep_chan_data_3_12 = out_chan_dep_data_3;
    assign token_3_12 = token_out_vec_3[12];
    assign dep_chan_vld_3_13 = out_chan_dep_vld_vec_3[13];
    assign dep_chan_data_3_13 = out_chan_dep_data_3;
    assign token_3_13 = token_out_vec_3[13];
    assign dep_chan_vld_3_14 = out_chan_dep_vld_vec_3[14];
    assign dep_chan_data_3_14 = out_chan_dep_data_3;
    assign token_3_14 = token_out_vec_3[14];
    assign dep_chan_vld_3_15 = out_chan_dep_vld_vec_3[15];
    assign dep_chan_data_3_15 = out_chan_dep_data_3;
    assign token_3_15 = token_out_vec_3[15];
    assign dep_chan_vld_3_16 = out_chan_dep_vld_vec_3[16];
    assign dep_chan_data_3_16 = out_chan_dep_data_3;
    assign token_3_16 = token_out_vec_3[16];
    assign dep_chan_vld_3_17 = out_chan_dep_vld_vec_3[17];
    assign dep_chan_data_3_17 = out_chan_dep_data_3;
    assign token_3_17 = token_out_vec_3[17];
    assign dep_chan_vld_3_18 = out_chan_dep_vld_vec_3[18];
    assign dep_chan_data_3_18 = out_chan_dep_data_3;
    assign token_3_18 = token_out_vec_3[18];

    // Process: load_value33_U0
    kernel_pr_hls_deadlock_detect_unit #(35, 4, 19, 19) kernel_pr_hls_deadlock_detect_unit_4 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_4),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_4),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_4),
        .token_in_vec(token_in_vec_4),
        .dl_detect_in(dl_detect_out),
        .origin(origin[4]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_4),
        .out_chan_dep_data(out_chan_dep_data_4),
        .token_out_vec(token_out_vec_4),
        .dl_detect_out(dl_in_vec[4]));

    assign proc_4_data_FIFO_blk[0] = 1'b0 | (~load_value33_U0.value_r_blk_n);
    assign proc_4_data_PIPO_blk[0] = 1'b0;
    assign proc_4_start_FIFO_blk[0] = 1'b0;
    assign proc_4_TLF_FIFO_blk[0] = 1'b0;
    assign proc_4_input_sync_blk[0] = 1'b0 | (ap_sync_load_value33_U0_ap_ready & load_value33_U0.ap_idle & ~ap_sync_kernel_pr_entry98_U0_ap_ready);
    assign proc_4_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_4[0] = dl_detect_out ? proc_dep_vld_vec_4_reg[0] : (proc_4_data_FIFO_blk[0] | proc_4_data_PIPO_blk[0] | proc_4_start_FIFO_blk[0] | proc_4_TLF_FIFO_blk[0] | proc_4_input_sync_blk[0] | proc_4_output_sync_blk[0]);
    assign proc_4_data_FIFO_blk[1] = 1'b0 | (~load_value33_U0.bipedge_size_blk_n) | (~load_value33_U0.bipedge_stream_V_V1_blk_n);
    assign proc_4_data_PIPO_blk[1] = 1'b0;
    assign proc_4_start_FIFO_blk[1] = 1'b0;
    assign proc_4_TLF_FIFO_blk[1] = 1'b0;
    assign proc_4_input_sync_blk[1] = 1'b0 | (ap_sync_load_value33_U0_ap_ready & load_value33_U0.ap_idle & ~ap_sync_load_bipedge30_U0_ap_ready);
    assign proc_4_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_4[1] = dl_detect_out ? proc_dep_vld_vec_4_reg[1] : (proc_4_data_FIFO_blk[1] | proc_4_data_PIPO_blk[1] | proc_4_start_FIFO_blk[1] | proc_4_TLF_FIFO_blk[1] | proc_4_input_sync_blk[1] | proc_4_output_sync_blk[1]);
    assign proc_4_data_FIFO_blk[2] = 1'b0 | (~load_value33_U0.value_stream_V_V16_blk_n);
    assign proc_4_data_PIPO_blk[2] = 1'b0;
    assign proc_4_start_FIFO_blk[2] = 1'b0;
    assign proc_4_TLF_FIFO_blk[2] = 1'b0;
    assign proc_4_input_sync_blk[2] = 1'b0;
    assign proc_4_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_4[2] = dl_detect_out ? proc_dep_vld_vec_4_reg[2] : (proc_4_data_FIFO_blk[2] | proc_4_data_PIPO_blk[2] | proc_4_start_FIFO_blk[2] | proc_4_TLF_FIFO_blk[2] | proc_4_input_sync_blk[2] | proc_4_output_sync_blk[2]);
    assign proc_4_data_FIFO_blk[3] = 1'b0;
    assign proc_4_data_PIPO_blk[3] = 1'b0;
    assign proc_4_start_FIFO_blk[3] = 1'b0;
    assign proc_4_TLF_FIFO_blk[3] = 1'b0;
    assign proc_4_input_sync_blk[3] = 1'b0 | (ap_sync_load_value33_U0_ap_ready & load_value33_U0.ap_idle & ~ap_sync_load_bipedge31_U0_ap_ready);
    assign proc_4_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_4[3] = dl_detect_out ? proc_dep_vld_vec_4_reg[3] : (proc_4_data_FIFO_blk[3] | proc_4_data_PIPO_blk[3] | proc_4_start_FIFO_blk[3] | proc_4_TLF_FIFO_blk[3] | proc_4_input_sync_blk[3] | proc_4_output_sync_blk[3]);
    assign proc_4_data_FIFO_blk[4] = 1'b0;
    assign proc_4_data_PIPO_blk[4] = 1'b0;
    assign proc_4_start_FIFO_blk[4] = 1'b0;
    assign proc_4_TLF_FIFO_blk[4] = 1'b0;
    assign proc_4_input_sync_blk[4] = 1'b0 | (ap_sync_load_value33_U0_ap_ready & load_value33_U0.ap_idle & ~ap_sync_load_value32_U0_ap_ready);
    assign proc_4_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_4[4] = dl_detect_out ? proc_dep_vld_vec_4_reg[4] : (proc_4_data_FIFO_blk[4] | proc_4_data_PIPO_blk[4] | proc_4_start_FIFO_blk[4] | proc_4_TLF_FIFO_blk[4] | proc_4_input_sync_blk[4] | proc_4_output_sync_blk[4]);
    assign proc_4_data_FIFO_blk[5] = 1'b0;
    assign proc_4_data_PIPO_blk[5] = 1'b0;
    assign proc_4_start_FIFO_blk[5] = 1'b0;
    assign proc_4_TLF_FIFO_blk[5] = 1'b0;
    assign proc_4_input_sync_blk[5] = 1'b0 | (ap_sync_load_value33_U0_ap_ready & load_value33_U0.ap_idle & ~ap_sync_load_value34_U0_ap_ready);
    assign proc_4_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_4[5] = dl_detect_out ? proc_dep_vld_vec_4_reg[5] : (proc_4_data_FIFO_blk[5] | proc_4_data_PIPO_blk[5] | proc_4_start_FIFO_blk[5] | proc_4_TLF_FIFO_blk[5] | proc_4_input_sync_blk[5] | proc_4_output_sync_blk[5]);
    assign proc_4_data_FIFO_blk[6] = 1'b0;
    assign proc_4_data_PIPO_blk[6] = 1'b0;
    assign proc_4_start_FIFO_blk[6] = 1'b0;
    assign proc_4_TLF_FIFO_blk[6] = 1'b0;
    assign proc_4_input_sync_blk[6] = 1'b0 | (ap_sync_load_value33_U0_ap_ready & load_value33_U0.ap_idle & ~ap_sync_load_value35_U0_ap_ready);
    assign proc_4_output_sync_blk[6] = 1'b0;
    assign proc_dep_vld_vec_4[6] = dl_detect_out ? proc_dep_vld_vec_4_reg[6] : (proc_4_data_FIFO_blk[6] | proc_4_data_PIPO_blk[6] | proc_4_start_FIFO_blk[6] | proc_4_TLF_FIFO_blk[6] | proc_4_input_sync_blk[6] | proc_4_output_sync_blk[6]);
    assign proc_4_data_FIFO_blk[7] = 1'b0;
    assign proc_4_data_PIPO_blk[7] = 1'b0;
    assign proc_4_start_FIFO_blk[7] = 1'b0;
    assign proc_4_TLF_FIFO_blk[7] = 1'b0;
    assign proc_4_input_sync_blk[7] = 1'b0 | (ap_sync_load_value33_U0_ap_ready & load_value33_U0.ap_idle & ~ap_sync_load_value36_U0_ap_ready);
    assign proc_4_output_sync_blk[7] = 1'b0;
    assign proc_dep_vld_vec_4[7] = dl_detect_out ? proc_dep_vld_vec_4_reg[7] : (proc_4_data_FIFO_blk[7] | proc_4_data_PIPO_blk[7] | proc_4_start_FIFO_blk[7] | proc_4_TLF_FIFO_blk[7] | proc_4_input_sync_blk[7] | proc_4_output_sync_blk[7]);
    assign proc_4_data_FIFO_blk[8] = 1'b0;
    assign proc_4_data_PIPO_blk[8] = 1'b0;
    assign proc_4_start_FIFO_blk[8] = 1'b0;
    assign proc_4_TLF_FIFO_blk[8] = 1'b0;
    assign proc_4_input_sync_blk[8] = 1'b0 | (ap_sync_load_value33_U0_ap_ready & load_value33_U0.ap_idle & ~ap_sync_load_value37_U0_ap_ready);
    assign proc_4_output_sync_blk[8] = 1'b0;
    assign proc_dep_vld_vec_4[8] = dl_detect_out ? proc_dep_vld_vec_4_reg[8] : (proc_4_data_FIFO_blk[8] | proc_4_data_PIPO_blk[8] | proc_4_start_FIFO_blk[8] | proc_4_TLF_FIFO_blk[8] | proc_4_input_sync_blk[8] | proc_4_output_sync_blk[8]);
    assign proc_4_data_FIFO_blk[9] = 1'b0;
    assign proc_4_data_PIPO_blk[9] = 1'b0;
    assign proc_4_start_FIFO_blk[9] = 1'b0;
    assign proc_4_TLF_FIFO_blk[9] = 1'b0;
    assign proc_4_input_sync_blk[9] = 1'b0 | (ap_sync_load_value33_U0_ap_ready & load_value33_U0.ap_idle & ~ap_sync_load_value38_U0_ap_ready);
    assign proc_4_output_sync_blk[9] = 1'b0;
    assign proc_dep_vld_vec_4[9] = dl_detect_out ? proc_dep_vld_vec_4_reg[9] : (proc_4_data_FIFO_blk[9] | proc_4_data_PIPO_blk[9] | proc_4_start_FIFO_blk[9] | proc_4_TLF_FIFO_blk[9] | proc_4_input_sync_blk[9] | proc_4_output_sync_blk[9]);
    assign proc_4_data_FIFO_blk[10] = 1'b0;
    assign proc_4_data_PIPO_blk[10] = 1'b0;
    assign proc_4_start_FIFO_blk[10] = 1'b0;
    assign proc_4_TLF_FIFO_blk[10] = 1'b0;
    assign proc_4_input_sync_blk[10] = 1'b0 | (ap_sync_load_value33_U0_ap_ready & load_value33_U0.ap_idle & ~ap_sync_load_value39_U0_ap_ready);
    assign proc_4_output_sync_blk[10] = 1'b0;
    assign proc_dep_vld_vec_4[10] = dl_detect_out ? proc_dep_vld_vec_4_reg[10] : (proc_4_data_FIFO_blk[10] | proc_4_data_PIPO_blk[10] | proc_4_start_FIFO_blk[10] | proc_4_TLF_FIFO_blk[10] | proc_4_input_sync_blk[10] | proc_4_output_sync_blk[10]);
    assign proc_4_data_FIFO_blk[11] = 1'b0;
    assign proc_4_data_PIPO_blk[11] = 1'b0;
    assign proc_4_start_FIFO_blk[11] = 1'b0;
    assign proc_4_TLF_FIFO_blk[11] = 1'b0;
    assign proc_4_input_sync_blk[11] = 1'b0 | (ap_sync_load_value33_U0_ap_ready & load_value33_U0.ap_idle & ~ap_sync_load_value40_U0_ap_ready);
    assign proc_4_output_sync_blk[11] = 1'b0;
    assign proc_dep_vld_vec_4[11] = dl_detect_out ? proc_dep_vld_vec_4_reg[11] : (proc_4_data_FIFO_blk[11] | proc_4_data_PIPO_blk[11] | proc_4_start_FIFO_blk[11] | proc_4_TLF_FIFO_blk[11] | proc_4_input_sync_blk[11] | proc_4_output_sync_blk[11]);
    assign proc_4_data_FIFO_blk[12] = 1'b0;
    assign proc_4_data_PIPO_blk[12] = 1'b0;
    assign proc_4_start_FIFO_blk[12] = 1'b0;
    assign proc_4_TLF_FIFO_blk[12] = 1'b0;
    assign proc_4_input_sync_blk[12] = 1'b0 | (ap_sync_load_value33_U0_ap_ready & load_value33_U0.ap_idle & ~ap_sync_load_value41_U0_ap_ready);
    assign proc_4_output_sync_blk[12] = 1'b0;
    assign proc_dep_vld_vec_4[12] = dl_detect_out ? proc_dep_vld_vec_4_reg[12] : (proc_4_data_FIFO_blk[12] | proc_4_data_PIPO_blk[12] | proc_4_start_FIFO_blk[12] | proc_4_TLF_FIFO_blk[12] | proc_4_input_sync_blk[12] | proc_4_output_sync_blk[12]);
    assign proc_4_data_FIFO_blk[13] = 1'b0;
    assign proc_4_data_PIPO_blk[13] = 1'b0;
    assign proc_4_start_FIFO_blk[13] = 1'b0;
    assign proc_4_TLF_FIFO_blk[13] = 1'b0;
    assign proc_4_input_sync_blk[13] = 1'b0 | (ap_sync_load_value33_U0_ap_ready & load_value33_U0.ap_idle & ~ap_sync_load_value42_U0_ap_ready);
    assign proc_4_output_sync_blk[13] = 1'b0;
    assign proc_dep_vld_vec_4[13] = dl_detect_out ? proc_dep_vld_vec_4_reg[13] : (proc_4_data_FIFO_blk[13] | proc_4_data_PIPO_blk[13] | proc_4_start_FIFO_blk[13] | proc_4_TLF_FIFO_blk[13] | proc_4_input_sync_blk[13] | proc_4_output_sync_blk[13]);
    assign proc_4_data_FIFO_blk[14] = 1'b0;
    assign proc_4_data_PIPO_blk[14] = 1'b0;
    assign proc_4_start_FIFO_blk[14] = 1'b0;
    assign proc_4_TLF_FIFO_blk[14] = 1'b0;
    assign proc_4_input_sync_blk[14] = 1'b0 | (ap_sync_load_value33_U0_ap_ready & load_value33_U0.ap_idle & ~ap_sync_load_value43_U0_ap_ready);
    assign proc_4_output_sync_blk[14] = 1'b0;
    assign proc_dep_vld_vec_4[14] = dl_detect_out ? proc_dep_vld_vec_4_reg[14] : (proc_4_data_FIFO_blk[14] | proc_4_data_PIPO_blk[14] | proc_4_start_FIFO_blk[14] | proc_4_TLF_FIFO_blk[14] | proc_4_input_sync_blk[14] | proc_4_output_sync_blk[14]);
    assign proc_4_data_FIFO_blk[15] = 1'b0;
    assign proc_4_data_PIPO_blk[15] = 1'b0;
    assign proc_4_start_FIFO_blk[15] = 1'b0;
    assign proc_4_TLF_FIFO_blk[15] = 1'b0;
    assign proc_4_input_sync_blk[15] = 1'b0 | (ap_sync_load_value33_U0_ap_ready & load_value33_U0.ap_idle & ~ap_sync_load_value44_U0_ap_ready);
    assign proc_4_output_sync_blk[15] = 1'b0;
    assign proc_dep_vld_vec_4[15] = dl_detect_out ? proc_dep_vld_vec_4_reg[15] : (proc_4_data_FIFO_blk[15] | proc_4_data_PIPO_blk[15] | proc_4_start_FIFO_blk[15] | proc_4_TLF_FIFO_blk[15] | proc_4_input_sync_blk[15] | proc_4_output_sync_blk[15]);
    assign proc_4_data_FIFO_blk[16] = 1'b0;
    assign proc_4_data_PIPO_blk[16] = 1'b0;
    assign proc_4_start_FIFO_blk[16] = 1'b0;
    assign proc_4_TLF_FIFO_blk[16] = 1'b0;
    assign proc_4_input_sync_blk[16] = 1'b0 | (ap_sync_load_value33_U0_ap_ready & load_value33_U0.ap_idle & ~ap_sync_load_value45_U0_ap_ready);
    assign proc_4_output_sync_blk[16] = 1'b0;
    assign proc_dep_vld_vec_4[16] = dl_detect_out ? proc_dep_vld_vec_4_reg[16] : (proc_4_data_FIFO_blk[16] | proc_4_data_PIPO_blk[16] | proc_4_start_FIFO_blk[16] | proc_4_TLF_FIFO_blk[16] | proc_4_input_sync_blk[16] | proc_4_output_sync_blk[16]);
    assign proc_4_data_FIFO_blk[17] = 1'b0;
    assign proc_4_data_PIPO_blk[17] = 1'b0;
    assign proc_4_start_FIFO_blk[17] = 1'b0;
    assign proc_4_TLF_FIFO_blk[17] = 1'b0;
    assign proc_4_input_sync_blk[17] = 1'b0 | (ap_sync_load_value33_U0_ap_ready & load_value33_U0.ap_idle & ~ap_sync_load_value46_U0_ap_ready);
    assign proc_4_output_sync_blk[17] = 1'b0;
    assign proc_dep_vld_vec_4[17] = dl_detect_out ? proc_dep_vld_vec_4_reg[17] : (proc_4_data_FIFO_blk[17] | proc_4_data_PIPO_blk[17] | proc_4_start_FIFO_blk[17] | proc_4_TLF_FIFO_blk[17] | proc_4_input_sync_blk[17] | proc_4_output_sync_blk[17]);
    assign proc_4_data_FIFO_blk[18] = 1'b0;
    assign proc_4_data_PIPO_blk[18] = 1'b0;
    assign proc_4_start_FIFO_blk[18] = 1'b0;
    assign proc_4_TLF_FIFO_blk[18] = 1'b0;
    assign proc_4_input_sync_blk[18] = 1'b0 | (ap_sync_load_value33_U0_ap_ready & load_value33_U0.ap_idle & ~ap_sync_load_value47_U0_ap_ready);
    assign proc_4_output_sync_blk[18] = 1'b0;
    assign proc_dep_vld_vec_4[18] = dl_detect_out ? proc_dep_vld_vec_4_reg[18] : (proc_4_data_FIFO_blk[18] | proc_4_data_PIPO_blk[18] | proc_4_start_FIFO_blk[18] | proc_4_TLF_FIFO_blk[18] | proc_4_input_sync_blk[18] | proc_4_output_sync_blk[18]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_4_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_4_reg <= proc_dep_vld_vec_4;
        end
    end
    assign in_chan_dep_vld_vec_4[0] = dep_chan_vld_0_4;
    assign in_chan_dep_data_vec_4[34 : 0] = dep_chan_data_0_4;
    assign token_in_vec_4[0] = token_0_4;
    assign in_chan_dep_vld_vec_4[1] = dep_chan_vld_1_4;
    assign in_chan_dep_data_vec_4[69 : 35] = dep_chan_data_1_4;
    assign token_in_vec_4[1] = token_1_4;
    assign in_chan_dep_vld_vec_4[2] = dep_chan_vld_2_4;
    assign in_chan_dep_data_vec_4[104 : 70] = dep_chan_data_2_4;
    assign token_in_vec_4[2] = token_2_4;
    assign in_chan_dep_vld_vec_4[3] = dep_chan_vld_3_4;
    assign in_chan_dep_data_vec_4[139 : 105] = dep_chan_data_3_4;
    assign token_in_vec_4[3] = token_3_4;
    assign in_chan_dep_vld_vec_4[4] = dep_chan_vld_5_4;
    assign in_chan_dep_data_vec_4[174 : 140] = dep_chan_data_5_4;
    assign token_in_vec_4[4] = token_5_4;
    assign in_chan_dep_vld_vec_4[5] = dep_chan_vld_6_4;
    assign in_chan_dep_data_vec_4[209 : 175] = dep_chan_data_6_4;
    assign token_in_vec_4[5] = token_6_4;
    assign in_chan_dep_vld_vec_4[6] = dep_chan_vld_7_4;
    assign in_chan_dep_data_vec_4[244 : 210] = dep_chan_data_7_4;
    assign token_in_vec_4[6] = token_7_4;
    assign in_chan_dep_vld_vec_4[7] = dep_chan_vld_8_4;
    assign in_chan_dep_data_vec_4[279 : 245] = dep_chan_data_8_4;
    assign token_in_vec_4[7] = token_8_4;
    assign in_chan_dep_vld_vec_4[8] = dep_chan_vld_9_4;
    assign in_chan_dep_data_vec_4[314 : 280] = dep_chan_data_9_4;
    assign token_in_vec_4[8] = token_9_4;
    assign in_chan_dep_vld_vec_4[9] = dep_chan_vld_10_4;
    assign in_chan_dep_data_vec_4[349 : 315] = dep_chan_data_10_4;
    assign token_in_vec_4[9] = token_10_4;
    assign in_chan_dep_vld_vec_4[10] = dep_chan_vld_11_4;
    assign in_chan_dep_data_vec_4[384 : 350] = dep_chan_data_11_4;
    assign token_in_vec_4[10] = token_11_4;
    assign in_chan_dep_vld_vec_4[11] = dep_chan_vld_12_4;
    assign in_chan_dep_data_vec_4[419 : 385] = dep_chan_data_12_4;
    assign token_in_vec_4[11] = token_12_4;
    assign in_chan_dep_vld_vec_4[12] = dep_chan_vld_13_4;
    assign in_chan_dep_data_vec_4[454 : 420] = dep_chan_data_13_4;
    assign token_in_vec_4[12] = token_13_4;
    assign in_chan_dep_vld_vec_4[13] = dep_chan_vld_14_4;
    assign in_chan_dep_data_vec_4[489 : 455] = dep_chan_data_14_4;
    assign token_in_vec_4[13] = token_14_4;
    assign in_chan_dep_vld_vec_4[14] = dep_chan_vld_15_4;
    assign in_chan_dep_data_vec_4[524 : 490] = dep_chan_data_15_4;
    assign token_in_vec_4[14] = token_15_4;
    assign in_chan_dep_vld_vec_4[15] = dep_chan_vld_16_4;
    assign in_chan_dep_data_vec_4[559 : 525] = dep_chan_data_16_4;
    assign token_in_vec_4[15] = token_16_4;
    assign in_chan_dep_vld_vec_4[16] = dep_chan_vld_17_4;
    assign in_chan_dep_data_vec_4[594 : 560] = dep_chan_data_17_4;
    assign token_in_vec_4[16] = token_17_4;
    assign in_chan_dep_vld_vec_4[17] = dep_chan_vld_18_4;
    assign in_chan_dep_data_vec_4[629 : 595] = dep_chan_data_18_4;
    assign token_in_vec_4[17] = token_18_4;
    assign in_chan_dep_vld_vec_4[18] = dep_chan_vld_20_4;
    assign in_chan_dep_data_vec_4[664 : 630] = dep_chan_data_20_4;
    assign token_in_vec_4[18] = token_20_4;
    assign dep_chan_vld_4_0 = out_chan_dep_vld_vec_4[0];
    assign dep_chan_data_4_0 = out_chan_dep_data_4;
    assign token_4_0 = token_out_vec_4[0];
    assign dep_chan_vld_4_1 = out_chan_dep_vld_vec_4[1];
    assign dep_chan_data_4_1 = out_chan_dep_data_4;
    assign token_4_1 = token_out_vec_4[1];
    assign dep_chan_vld_4_20 = out_chan_dep_vld_vec_4[2];
    assign dep_chan_data_4_20 = out_chan_dep_data_4;
    assign token_4_20 = token_out_vec_4[2];
    assign dep_chan_vld_4_2 = out_chan_dep_vld_vec_4[3];
    assign dep_chan_data_4_2 = out_chan_dep_data_4;
    assign token_4_2 = token_out_vec_4[3];
    assign dep_chan_vld_4_3 = out_chan_dep_vld_vec_4[4];
    assign dep_chan_data_4_3 = out_chan_dep_data_4;
    assign token_4_3 = token_out_vec_4[4];
    assign dep_chan_vld_4_5 = out_chan_dep_vld_vec_4[5];
    assign dep_chan_data_4_5 = out_chan_dep_data_4;
    assign token_4_5 = token_out_vec_4[5];
    assign dep_chan_vld_4_6 = out_chan_dep_vld_vec_4[6];
    assign dep_chan_data_4_6 = out_chan_dep_data_4;
    assign token_4_6 = token_out_vec_4[6];
    assign dep_chan_vld_4_7 = out_chan_dep_vld_vec_4[7];
    assign dep_chan_data_4_7 = out_chan_dep_data_4;
    assign token_4_7 = token_out_vec_4[7];
    assign dep_chan_vld_4_8 = out_chan_dep_vld_vec_4[8];
    assign dep_chan_data_4_8 = out_chan_dep_data_4;
    assign token_4_8 = token_out_vec_4[8];
    assign dep_chan_vld_4_9 = out_chan_dep_vld_vec_4[9];
    assign dep_chan_data_4_9 = out_chan_dep_data_4;
    assign token_4_9 = token_out_vec_4[9];
    assign dep_chan_vld_4_10 = out_chan_dep_vld_vec_4[10];
    assign dep_chan_data_4_10 = out_chan_dep_data_4;
    assign token_4_10 = token_out_vec_4[10];
    assign dep_chan_vld_4_11 = out_chan_dep_vld_vec_4[11];
    assign dep_chan_data_4_11 = out_chan_dep_data_4;
    assign token_4_11 = token_out_vec_4[11];
    assign dep_chan_vld_4_12 = out_chan_dep_vld_vec_4[12];
    assign dep_chan_data_4_12 = out_chan_dep_data_4;
    assign token_4_12 = token_out_vec_4[12];
    assign dep_chan_vld_4_13 = out_chan_dep_vld_vec_4[13];
    assign dep_chan_data_4_13 = out_chan_dep_data_4;
    assign token_4_13 = token_out_vec_4[13];
    assign dep_chan_vld_4_14 = out_chan_dep_vld_vec_4[14];
    assign dep_chan_data_4_14 = out_chan_dep_data_4;
    assign token_4_14 = token_out_vec_4[14];
    assign dep_chan_vld_4_15 = out_chan_dep_vld_vec_4[15];
    assign dep_chan_data_4_15 = out_chan_dep_data_4;
    assign token_4_15 = token_out_vec_4[15];
    assign dep_chan_vld_4_16 = out_chan_dep_vld_vec_4[16];
    assign dep_chan_data_4_16 = out_chan_dep_data_4;
    assign token_4_16 = token_out_vec_4[16];
    assign dep_chan_vld_4_17 = out_chan_dep_vld_vec_4[17];
    assign dep_chan_data_4_17 = out_chan_dep_data_4;
    assign token_4_17 = token_out_vec_4[17];
    assign dep_chan_vld_4_18 = out_chan_dep_vld_vec_4[18];
    assign dep_chan_data_4_18 = out_chan_dep_data_4;
    assign token_4_18 = token_out_vec_4[18];

    // Process: load_value34_U0
    kernel_pr_hls_deadlock_detect_unit #(35, 5, 19, 19) kernel_pr_hls_deadlock_detect_unit_5 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_5),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_5),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_5),
        .token_in_vec(token_in_vec_5),
        .dl_detect_in(dl_detect_out),
        .origin(origin[5]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_5),
        .out_chan_dep_data(out_chan_dep_data_5),
        .token_out_vec(token_out_vec_5),
        .dl_detect_out(dl_in_vec[5]));

    assign proc_5_data_FIFO_blk[0] = 1'b0 | (~load_value34_U0.value_r_blk_n);
    assign proc_5_data_PIPO_blk[0] = 1'b0;
    assign proc_5_start_FIFO_blk[0] = 1'b0;
    assign proc_5_TLF_FIFO_blk[0] = 1'b0;
    assign proc_5_input_sync_blk[0] = 1'b0 | (ap_sync_load_value34_U0_ap_ready & load_value34_U0.ap_idle & ~ap_sync_kernel_pr_entry98_U0_ap_ready);
    assign proc_5_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_5[0] = dl_detect_out ? proc_dep_vld_vec_5_reg[0] : (proc_5_data_FIFO_blk[0] | proc_5_data_PIPO_blk[0] | proc_5_start_FIFO_blk[0] | proc_5_TLF_FIFO_blk[0] | proc_5_input_sync_blk[0] | proc_5_output_sync_blk[0]);
    assign proc_5_data_FIFO_blk[1] = 1'b0 | (~load_value34_U0.bipedge_size_blk_n) | (~load_value34_U0.bipedge_stream_V_V2_blk_n);
    assign proc_5_data_PIPO_blk[1] = 1'b0;
    assign proc_5_start_FIFO_blk[1] = 1'b0;
    assign proc_5_TLF_FIFO_blk[1] = 1'b0;
    assign proc_5_input_sync_blk[1] = 1'b0 | (ap_sync_load_value34_U0_ap_ready & load_value34_U0.ap_idle & ~ap_sync_load_bipedge30_U0_ap_ready);
    assign proc_5_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_5[1] = dl_detect_out ? proc_dep_vld_vec_5_reg[1] : (proc_5_data_FIFO_blk[1] | proc_5_data_PIPO_blk[1] | proc_5_start_FIFO_blk[1] | proc_5_TLF_FIFO_blk[1] | proc_5_input_sync_blk[1] | proc_5_output_sync_blk[1]);
    assign proc_5_data_FIFO_blk[2] = 1'b0 | (~load_value34_U0.value_stream_V_V17_blk_n);
    assign proc_5_data_PIPO_blk[2] = 1'b0;
    assign proc_5_start_FIFO_blk[2] = 1'b0;
    assign proc_5_TLF_FIFO_blk[2] = 1'b0;
    assign proc_5_input_sync_blk[2] = 1'b0;
    assign proc_5_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_5[2] = dl_detect_out ? proc_dep_vld_vec_5_reg[2] : (proc_5_data_FIFO_blk[2] | proc_5_data_PIPO_blk[2] | proc_5_start_FIFO_blk[2] | proc_5_TLF_FIFO_blk[2] | proc_5_input_sync_blk[2] | proc_5_output_sync_blk[2]);
    assign proc_5_data_FIFO_blk[3] = 1'b0;
    assign proc_5_data_PIPO_blk[3] = 1'b0;
    assign proc_5_start_FIFO_blk[3] = 1'b0;
    assign proc_5_TLF_FIFO_blk[3] = 1'b0;
    assign proc_5_input_sync_blk[3] = 1'b0 | (ap_sync_load_value34_U0_ap_ready & load_value34_U0.ap_idle & ~ap_sync_load_bipedge31_U0_ap_ready);
    assign proc_5_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_5[3] = dl_detect_out ? proc_dep_vld_vec_5_reg[3] : (proc_5_data_FIFO_blk[3] | proc_5_data_PIPO_blk[3] | proc_5_start_FIFO_blk[3] | proc_5_TLF_FIFO_blk[3] | proc_5_input_sync_blk[3] | proc_5_output_sync_blk[3]);
    assign proc_5_data_FIFO_blk[4] = 1'b0;
    assign proc_5_data_PIPO_blk[4] = 1'b0;
    assign proc_5_start_FIFO_blk[4] = 1'b0;
    assign proc_5_TLF_FIFO_blk[4] = 1'b0;
    assign proc_5_input_sync_blk[4] = 1'b0 | (ap_sync_load_value34_U0_ap_ready & load_value34_U0.ap_idle & ~ap_sync_load_value32_U0_ap_ready);
    assign proc_5_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_5[4] = dl_detect_out ? proc_dep_vld_vec_5_reg[4] : (proc_5_data_FIFO_blk[4] | proc_5_data_PIPO_blk[4] | proc_5_start_FIFO_blk[4] | proc_5_TLF_FIFO_blk[4] | proc_5_input_sync_blk[4] | proc_5_output_sync_blk[4]);
    assign proc_5_data_FIFO_blk[5] = 1'b0;
    assign proc_5_data_PIPO_blk[5] = 1'b0;
    assign proc_5_start_FIFO_blk[5] = 1'b0;
    assign proc_5_TLF_FIFO_blk[5] = 1'b0;
    assign proc_5_input_sync_blk[5] = 1'b0 | (ap_sync_load_value34_U0_ap_ready & load_value34_U0.ap_idle & ~ap_sync_load_value33_U0_ap_ready);
    assign proc_5_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_5[5] = dl_detect_out ? proc_dep_vld_vec_5_reg[5] : (proc_5_data_FIFO_blk[5] | proc_5_data_PIPO_blk[5] | proc_5_start_FIFO_blk[5] | proc_5_TLF_FIFO_blk[5] | proc_5_input_sync_blk[5] | proc_5_output_sync_blk[5]);
    assign proc_5_data_FIFO_blk[6] = 1'b0;
    assign proc_5_data_PIPO_blk[6] = 1'b0;
    assign proc_5_start_FIFO_blk[6] = 1'b0;
    assign proc_5_TLF_FIFO_blk[6] = 1'b0;
    assign proc_5_input_sync_blk[6] = 1'b0 | (ap_sync_load_value34_U0_ap_ready & load_value34_U0.ap_idle & ~ap_sync_load_value35_U0_ap_ready);
    assign proc_5_output_sync_blk[6] = 1'b0;
    assign proc_dep_vld_vec_5[6] = dl_detect_out ? proc_dep_vld_vec_5_reg[6] : (proc_5_data_FIFO_blk[6] | proc_5_data_PIPO_blk[6] | proc_5_start_FIFO_blk[6] | proc_5_TLF_FIFO_blk[6] | proc_5_input_sync_blk[6] | proc_5_output_sync_blk[6]);
    assign proc_5_data_FIFO_blk[7] = 1'b0;
    assign proc_5_data_PIPO_blk[7] = 1'b0;
    assign proc_5_start_FIFO_blk[7] = 1'b0;
    assign proc_5_TLF_FIFO_blk[7] = 1'b0;
    assign proc_5_input_sync_blk[7] = 1'b0 | (ap_sync_load_value34_U0_ap_ready & load_value34_U0.ap_idle & ~ap_sync_load_value36_U0_ap_ready);
    assign proc_5_output_sync_blk[7] = 1'b0;
    assign proc_dep_vld_vec_5[7] = dl_detect_out ? proc_dep_vld_vec_5_reg[7] : (proc_5_data_FIFO_blk[7] | proc_5_data_PIPO_blk[7] | proc_5_start_FIFO_blk[7] | proc_5_TLF_FIFO_blk[7] | proc_5_input_sync_blk[7] | proc_5_output_sync_blk[7]);
    assign proc_5_data_FIFO_blk[8] = 1'b0;
    assign proc_5_data_PIPO_blk[8] = 1'b0;
    assign proc_5_start_FIFO_blk[8] = 1'b0;
    assign proc_5_TLF_FIFO_blk[8] = 1'b0;
    assign proc_5_input_sync_blk[8] = 1'b0 | (ap_sync_load_value34_U0_ap_ready & load_value34_U0.ap_idle & ~ap_sync_load_value37_U0_ap_ready);
    assign proc_5_output_sync_blk[8] = 1'b0;
    assign proc_dep_vld_vec_5[8] = dl_detect_out ? proc_dep_vld_vec_5_reg[8] : (proc_5_data_FIFO_blk[8] | proc_5_data_PIPO_blk[8] | proc_5_start_FIFO_blk[8] | proc_5_TLF_FIFO_blk[8] | proc_5_input_sync_blk[8] | proc_5_output_sync_blk[8]);
    assign proc_5_data_FIFO_blk[9] = 1'b0;
    assign proc_5_data_PIPO_blk[9] = 1'b0;
    assign proc_5_start_FIFO_blk[9] = 1'b0;
    assign proc_5_TLF_FIFO_blk[9] = 1'b0;
    assign proc_5_input_sync_blk[9] = 1'b0 | (ap_sync_load_value34_U0_ap_ready & load_value34_U0.ap_idle & ~ap_sync_load_value38_U0_ap_ready);
    assign proc_5_output_sync_blk[9] = 1'b0;
    assign proc_dep_vld_vec_5[9] = dl_detect_out ? proc_dep_vld_vec_5_reg[9] : (proc_5_data_FIFO_blk[9] | proc_5_data_PIPO_blk[9] | proc_5_start_FIFO_blk[9] | proc_5_TLF_FIFO_blk[9] | proc_5_input_sync_blk[9] | proc_5_output_sync_blk[9]);
    assign proc_5_data_FIFO_blk[10] = 1'b0;
    assign proc_5_data_PIPO_blk[10] = 1'b0;
    assign proc_5_start_FIFO_blk[10] = 1'b0;
    assign proc_5_TLF_FIFO_blk[10] = 1'b0;
    assign proc_5_input_sync_blk[10] = 1'b0 | (ap_sync_load_value34_U0_ap_ready & load_value34_U0.ap_idle & ~ap_sync_load_value39_U0_ap_ready);
    assign proc_5_output_sync_blk[10] = 1'b0;
    assign proc_dep_vld_vec_5[10] = dl_detect_out ? proc_dep_vld_vec_5_reg[10] : (proc_5_data_FIFO_blk[10] | proc_5_data_PIPO_blk[10] | proc_5_start_FIFO_blk[10] | proc_5_TLF_FIFO_blk[10] | proc_5_input_sync_blk[10] | proc_5_output_sync_blk[10]);
    assign proc_5_data_FIFO_blk[11] = 1'b0;
    assign proc_5_data_PIPO_blk[11] = 1'b0;
    assign proc_5_start_FIFO_blk[11] = 1'b0;
    assign proc_5_TLF_FIFO_blk[11] = 1'b0;
    assign proc_5_input_sync_blk[11] = 1'b0 | (ap_sync_load_value34_U0_ap_ready & load_value34_U0.ap_idle & ~ap_sync_load_value40_U0_ap_ready);
    assign proc_5_output_sync_blk[11] = 1'b0;
    assign proc_dep_vld_vec_5[11] = dl_detect_out ? proc_dep_vld_vec_5_reg[11] : (proc_5_data_FIFO_blk[11] | proc_5_data_PIPO_blk[11] | proc_5_start_FIFO_blk[11] | proc_5_TLF_FIFO_blk[11] | proc_5_input_sync_blk[11] | proc_5_output_sync_blk[11]);
    assign proc_5_data_FIFO_blk[12] = 1'b0;
    assign proc_5_data_PIPO_blk[12] = 1'b0;
    assign proc_5_start_FIFO_blk[12] = 1'b0;
    assign proc_5_TLF_FIFO_blk[12] = 1'b0;
    assign proc_5_input_sync_blk[12] = 1'b0 | (ap_sync_load_value34_U0_ap_ready & load_value34_U0.ap_idle & ~ap_sync_load_value41_U0_ap_ready);
    assign proc_5_output_sync_blk[12] = 1'b0;
    assign proc_dep_vld_vec_5[12] = dl_detect_out ? proc_dep_vld_vec_5_reg[12] : (proc_5_data_FIFO_blk[12] | proc_5_data_PIPO_blk[12] | proc_5_start_FIFO_blk[12] | proc_5_TLF_FIFO_blk[12] | proc_5_input_sync_blk[12] | proc_5_output_sync_blk[12]);
    assign proc_5_data_FIFO_blk[13] = 1'b0;
    assign proc_5_data_PIPO_blk[13] = 1'b0;
    assign proc_5_start_FIFO_blk[13] = 1'b0;
    assign proc_5_TLF_FIFO_blk[13] = 1'b0;
    assign proc_5_input_sync_blk[13] = 1'b0 | (ap_sync_load_value34_U0_ap_ready & load_value34_U0.ap_idle & ~ap_sync_load_value42_U0_ap_ready);
    assign proc_5_output_sync_blk[13] = 1'b0;
    assign proc_dep_vld_vec_5[13] = dl_detect_out ? proc_dep_vld_vec_5_reg[13] : (proc_5_data_FIFO_blk[13] | proc_5_data_PIPO_blk[13] | proc_5_start_FIFO_blk[13] | proc_5_TLF_FIFO_blk[13] | proc_5_input_sync_blk[13] | proc_5_output_sync_blk[13]);
    assign proc_5_data_FIFO_blk[14] = 1'b0;
    assign proc_5_data_PIPO_blk[14] = 1'b0;
    assign proc_5_start_FIFO_blk[14] = 1'b0;
    assign proc_5_TLF_FIFO_blk[14] = 1'b0;
    assign proc_5_input_sync_blk[14] = 1'b0 | (ap_sync_load_value34_U0_ap_ready & load_value34_U0.ap_idle & ~ap_sync_load_value43_U0_ap_ready);
    assign proc_5_output_sync_blk[14] = 1'b0;
    assign proc_dep_vld_vec_5[14] = dl_detect_out ? proc_dep_vld_vec_5_reg[14] : (proc_5_data_FIFO_blk[14] | proc_5_data_PIPO_blk[14] | proc_5_start_FIFO_blk[14] | proc_5_TLF_FIFO_blk[14] | proc_5_input_sync_blk[14] | proc_5_output_sync_blk[14]);
    assign proc_5_data_FIFO_blk[15] = 1'b0;
    assign proc_5_data_PIPO_blk[15] = 1'b0;
    assign proc_5_start_FIFO_blk[15] = 1'b0;
    assign proc_5_TLF_FIFO_blk[15] = 1'b0;
    assign proc_5_input_sync_blk[15] = 1'b0 | (ap_sync_load_value34_U0_ap_ready & load_value34_U0.ap_idle & ~ap_sync_load_value44_U0_ap_ready);
    assign proc_5_output_sync_blk[15] = 1'b0;
    assign proc_dep_vld_vec_5[15] = dl_detect_out ? proc_dep_vld_vec_5_reg[15] : (proc_5_data_FIFO_blk[15] | proc_5_data_PIPO_blk[15] | proc_5_start_FIFO_blk[15] | proc_5_TLF_FIFO_blk[15] | proc_5_input_sync_blk[15] | proc_5_output_sync_blk[15]);
    assign proc_5_data_FIFO_blk[16] = 1'b0;
    assign proc_5_data_PIPO_blk[16] = 1'b0;
    assign proc_5_start_FIFO_blk[16] = 1'b0;
    assign proc_5_TLF_FIFO_blk[16] = 1'b0;
    assign proc_5_input_sync_blk[16] = 1'b0 | (ap_sync_load_value34_U0_ap_ready & load_value34_U0.ap_idle & ~ap_sync_load_value45_U0_ap_ready);
    assign proc_5_output_sync_blk[16] = 1'b0;
    assign proc_dep_vld_vec_5[16] = dl_detect_out ? proc_dep_vld_vec_5_reg[16] : (proc_5_data_FIFO_blk[16] | proc_5_data_PIPO_blk[16] | proc_5_start_FIFO_blk[16] | proc_5_TLF_FIFO_blk[16] | proc_5_input_sync_blk[16] | proc_5_output_sync_blk[16]);
    assign proc_5_data_FIFO_blk[17] = 1'b0;
    assign proc_5_data_PIPO_blk[17] = 1'b0;
    assign proc_5_start_FIFO_blk[17] = 1'b0;
    assign proc_5_TLF_FIFO_blk[17] = 1'b0;
    assign proc_5_input_sync_blk[17] = 1'b0 | (ap_sync_load_value34_U0_ap_ready & load_value34_U0.ap_idle & ~ap_sync_load_value46_U0_ap_ready);
    assign proc_5_output_sync_blk[17] = 1'b0;
    assign proc_dep_vld_vec_5[17] = dl_detect_out ? proc_dep_vld_vec_5_reg[17] : (proc_5_data_FIFO_blk[17] | proc_5_data_PIPO_blk[17] | proc_5_start_FIFO_blk[17] | proc_5_TLF_FIFO_blk[17] | proc_5_input_sync_blk[17] | proc_5_output_sync_blk[17]);
    assign proc_5_data_FIFO_blk[18] = 1'b0;
    assign proc_5_data_PIPO_blk[18] = 1'b0;
    assign proc_5_start_FIFO_blk[18] = 1'b0;
    assign proc_5_TLF_FIFO_blk[18] = 1'b0;
    assign proc_5_input_sync_blk[18] = 1'b0 | (ap_sync_load_value34_U0_ap_ready & load_value34_U0.ap_idle & ~ap_sync_load_value47_U0_ap_ready);
    assign proc_5_output_sync_blk[18] = 1'b0;
    assign proc_dep_vld_vec_5[18] = dl_detect_out ? proc_dep_vld_vec_5_reg[18] : (proc_5_data_FIFO_blk[18] | proc_5_data_PIPO_blk[18] | proc_5_start_FIFO_blk[18] | proc_5_TLF_FIFO_blk[18] | proc_5_input_sync_blk[18] | proc_5_output_sync_blk[18]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_5_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_5_reg <= proc_dep_vld_vec_5;
        end
    end
    assign in_chan_dep_vld_vec_5[0] = dep_chan_vld_0_5;
    assign in_chan_dep_data_vec_5[34 : 0] = dep_chan_data_0_5;
    assign token_in_vec_5[0] = token_0_5;
    assign in_chan_dep_vld_vec_5[1] = dep_chan_vld_1_5;
    assign in_chan_dep_data_vec_5[69 : 35] = dep_chan_data_1_5;
    assign token_in_vec_5[1] = token_1_5;
    assign in_chan_dep_vld_vec_5[2] = dep_chan_vld_2_5;
    assign in_chan_dep_data_vec_5[104 : 70] = dep_chan_data_2_5;
    assign token_in_vec_5[2] = token_2_5;
    assign in_chan_dep_vld_vec_5[3] = dep_chan_vld_3_5;
    assign in_chan_dep_data_vec_5[139 : 105] = dep_chan_data_3_5;
    assign token_in_vec_5[3] = token_3_5;
    assign in_chan_dep_vld_vec_5[4] = dep_chan_vld_4_5;
    assign in_chan_dep_data_vec_5[174 : 140] = dep_chan_data_4_5;
    assign token_in_vec_5[4] = token_4_5;
    assign in_chan_dep_vld_vec_5[5] = dep_chan_vld_6_5;
    assign in_chan_dep_data_vec_5[209 : 175] = dep_chan_data_6_5;
    assign token_in_vec_5[5] = token_6_5;
    assign in_chan_dep_vld_vec_5[6] = dep_chan_vld_7_5;
    assign in_chan_dep_data_vec_5[244 : 210] = dep_chan_data_7_5;
    assign token_in_vec_5[6] = token_7_5;
    assign in_chan_dep_vld_vec_5[7] = dep_chan_vld_8_5;
    assign in_chan_dep_data_vec_5[279 : 245] = dep_chan_data_8_5;
    assign token_in_vec_5[7] = token_8_5;
    assign in_chan_dep_vld_vec_5[8] = dep_chan_vld_9_5;
    assign in_chan_dep_data_vec_5[314 : 280] = dep_chan_data_9_5;
    assign token_in_vec_5[8] = token_9_5;
    assign in_chan_dep_vld_vec_5[9] = dep_chan_vld_10_5;
    assign in_chan_dep_data_vec_5[349 : 315] = dep_chan_data_10_5;
    assign token_in_vec_5[9] = token_10_5;
    assign in_chan_dep_vld_vec_5[10] = dep_chan_vld_11_5;
    assign in_chan_dep_data_vec_5[384 : 350] = dep_chan_data_11_5;
    assign token_in_vec_5[10] = token_11_5;
    assign in_chan_dep_vld_vec_5[11] = dep_chan_vld_12_5;
    assign in_chan_dep_data_vec_5[419 : 385] = dep_chan_data_12_5;
    assign token_in_vec_5[11] = token_12_5;
    assign in_chan_dep_vld_vec_5[12] = dep_chan_vld_13_5;
    assign in_chan_dep_data_vec_5[454 : 420] = dep_chan_data_13_5;
    assign token_in_vec_5[12] = token_13_5;
    assign in_chan_dep_vld_vec_5[13] = dep_chan_vld_14_5;
    assign in_chan_dep_data_vec_5[489 : 455] = dep_chan_data_14_5;
    assign token_in_vec_5[13] = token_14_5;
    assign in_chan_dep_vld_vec_5[14] = dep_chan_vld_15_5;
    assign in_chan_dep_data_vec_5[524 : 490] = dep_chan_data_15_5;
    assign token_in_vec_5[14] = token_15_5;
    assign in_chan_dep_vld_vec_5[15] = dep_chan_vld_16_5;
    assign in_chan_dep_data_vec_5[559 : 525] = dep_chan_data_16_5;
    assign token_in_vec_5[15] = token_16_5;
    assign in_chan_dep_vld_vec_5[16] = dep_chan_vld_17_5;
    assign in_chan_dep_data_vec_5[594 : 560] = dep_chan_data_17_5;
    assign token_in_vec_5[16] = token_17_5;
    assign in_chan_dep_vld_vec_5[17] = dep_chan_vld_18_5;
    assign in_chan_dep_data_vec_5[629 : 595] = dep_chan_data_18_5;
    assign token_in_vec_5[17] = token_18_5;
    assign in_chan_dep_vld_vec_5[18] = dep_chan_vld_21_5;
    assign in_chan_dep_data_vec_5[664 : 630] = dep_chan_data_21_5;
    assign token_in_vec_5[18] = token_21_5;
    assign dep_chan_vld_5_0 = out_chan_dep_vld_vec_5[0];
    assign dep_chan_data_5_0 = out_chan_dep_data_5;
    assign token_5_0 = token_out_vec_5[0];
    assign dep_chan_vld_5_1 = out_chan_dep_vld_vec_5[1];
    assign dep_chan_data_5_1 = out_chan_dep_data_5;
    assign token_5_1 = token_out_vec_5[1];
    assign dep_chan_vld_5_21 = out_chan_dep_vld_vec_5[2];
    assign dep_chan_data_5_21 = out_chan_dep_data_5;
    assign token_5_21 = token_out_vec_5[2];
    assign dep_chan_vld_5_2 = out_chan_dep_vld_vec_5[3];
    assign dep_chan_data_5_2 = out_chan_dep_data_5;
    assign token_5_2 = token_out_vec_5[3];
    assign dep_chan_vld_5_3 = out_chan_dep_vld_vec_5[4];
    assign dep_chan_data_5_3 = out_chan_dep_data_5;
    assign token_5_3 = token_out_vec_5[4];
    assign dep_chan_vld_5_4 = out_chan_dep_vld_vec_5[5];
    assign dep_chan_data_5_4 = out_chan_dep_data_5;
    assign token_5_4 = token_out_vec_5[5];
    assign dep_chan_vld_5_6 = out_chan_dep_vld_vec_5[6];
    assign dep_chan_data_5_6 = out_chan_dep_data_5;
    assign token_5_6 = token_out_vec_5[6];
    assign dep_chan_vld_5_7 = out_chan_dep_vld_vec_5[7];
    assign dep_chan_data_5_7 = out_chan_dep_data_5;
    assign token_5_7 = token_out_vec_5[7];
    assign dep_chan_vld_5_8 = out_chan_dep_vld_vec_5[8];
    assign dep_chan_data_5_8 = out_chan_dep_data_5;
    assign token_5_8 = token_out_vec_5[8];
    assign dep_chan_vld_5_9 = out_chan_dep_vld_vec_5[9];
    assign dep_chan_data_5_9 = out_chan_dep_data_5;
    assign token_5_9 = token_out_vec_5[9];
    assign dep_chan_vld_5_10 = out_chan_dep_vld_vec_5[10];
    assign dep_chan_data_5_10 = out_chan_dep_data_5;
    assign token_5_10 = token_out_vec_5[10];
    assign dep_chan_vld_5_11 = out_chan_dep_vld_vec_5[11];
    assign dep_chan_data_5_11 = out_chan_dep_data_5;
    assign token_5_11 = token_out_vec_5[11];
    assign dep_chan_vld_5_12 = out_chan_dep_vld_vec_5[12];
    assign dep_chan_data_5_12 = out_chan_dep_data_5;
    assign token_5_12 = token_out_vec_5[12];
    assign dep_chan_vld_5_13 = out_chan_dep_vld_vec_5[13];
    assign dep_chan_data_5_13 = out_chan_dep_data_5;
    assign token_5_13 = token_out_vec_5[13];
    assign dep_chan_vld_5_14 = out_chan_dep_vld_vec_5[14];
    assign dep_chan_data_5_14 = out_chan_dep_data_5;
    assign token_5_14 = token_out_vec_5[14];
    assign dep_chan_vld_5_15 = out_chan_dep_vld_vec_5[15];
    assign dep_chan_data_5_15 = out_chan_dep_data_5;
    assign token_5_15 = token_out_vec_5[15];
    assign dep_chan_vld_5_16 = out_chan_dep_vld_vec_5[16];
    assign dep_chan_data_5_16 = out_chan_dep_data_5;
    assign token_5_16 = token_out_vec_5[16];
    assign dep_chan_vld_5_17 = out_chan_dep_vld_vec_5[17];
    assign dep_chan_data_5_17 = out_chan_dep_data_5;
    assign token_5_17 = token_out_vec_5[17];
    assign dep_chan_vld_5_18 = out_chan_dep_vld_vec_5[18];
    assign dep_chan_data_5_18 = out_chan_dep_data_5;
    assign token_5_18 = token_out_vec_5[18];

    // Process: load_value35_U0
    kernel_pr_hls_deadlock_detect_unit #(35, 6, 19, 19) kernel_pr_hls_deadlock_detect_unit_6 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_6),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_6),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_6),
        .token_in_vec(token_in_vec_6),
        .dl_detect_in(dl_detect_out),
        .origin(origin[6]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_6),
        .out_chan_dep_data(out_chan_dep_data_6),
        .token_out_vec(token_out_vec_6),
        .dl_detect_out(dl_in_vec[6]));

    assign proc_6_data_FIFO_blk[0] = 1'b0 | (~load_value35_U0.value_r_blk_n);
    assign proc_6_data_PIPO_blk[0] = 1'b0;
    assign proc_6_start_FIFO_blk[0] = 1'b0;
    assign proc_6_TLF_FIFO_blk[0] = 1'b0;
    assign proc_6_input_sync_blk[0] = 1'b0 | (ap_sync_load_value35_U0_ap_ready & load_value35_U0.ap_idle & ~ap_sync_kernel_pr_entry98_U0_ap_ready);
    assign proc_6_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_6[0] = dl_detect_out ? proc_dep_vld_vec_6_reg[0] : (proc_6_data_FIFO_blk[0] | proc_6_data_PIPO_blk[0] | proc_6_start_FIFO_blk[0] | proc_6_TLF_FIFO_blk[0] | proc_6_input_sync_blk[0] | proc_6_output_sync_blk[0]);
    assign proc_6_data_FIFO_blk[1] = 1'b0 | (~load_value35_U0.bipedge_size_blk_n) | (~load_value35_U0.bipedge_stream_V_V3_blk_n);
    assign proc_6_data_PIPO_blk[1] = 1'b0;
    assign proc_6_start_FIFO_blk[1] = 1'b0;
    assign proc_6_TLF_FIFO_blk[1] = 1'b0;
    assign proc_6_input_sync_blk[1] = 1'b0 | (ap_sync_load_value35_U0_ap_ready & load_value35_U0.ap_idle & ~ap_sync_load_bipedge30_U0_ap_ready);
    assign proc_6_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_6[1] = dl_detect_out ? proc_dep_vld_vec_6_reg[1] : (proc_6_data_FIFO_blk[1] | proc_6_data_PIPO_blk[1] | proc_6_start_FIFO_blk[1] | proc_6_TLF_FIFO_blk[1] | proc_6_input_sync_blk[1] | proc_6_output_sync_blk[1]);
    assign proc_6_data_FIFO_blk[2] = 1'b0 | (~load_value35_U0.value_stream_V_V18_blk_n);
    assign proc_6_data_PIPO_blk[2] = 1'b0;
    assign proc_6_start_FIFO_blk[2] = 1'b0;
    assign proc_6_TLF_FIFO_blk[2] = 1'b0;
    assign proc_6_input_sync_blk[2] = 1'b0;
    assign proc_6_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_6[2] = dl_detect_out ? proc_dep_vld_vec_6_reg[2] : (proc_6_data_FIFO_blk[2] | proc_6_data_PIPO_blk[2] | proc_6_start_FIFO_blk[2] | proc_6_TLF_FIFO_blk[2] | proc_6_input_sync_blk[2] | proc_6_output_sync_blk[2]);
    assign proc_6_data_FIFO_blk[3] = 1'b0;
    assign proc_6_data_PIPO_blk[3] = 1'b0;
    assign proc_6_start_FIFO_blk[3] = 1'b0;
    assign proc_6_TLF_FIFO_blk[3] = 1'b0;
    assign proc_6_input_sync_blk[3] = 1'b0 | (ap_sync_load_value35_U0_ap_ready & load_value35_U0.ap_idle & ~ap_sync_load_bipedge31_U0_ap_ready);
    assign proc_6_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_6[3] = dl_detect_out ? proc_dep_vld_vec_6_reg[3] : (proc_6_data_FIFO_blk[3] | proc_6_data_PIPO_blk[3] | proc_6_start_FIFO_blk[3] | proc_6_TLF_FIFO_blk[3] | proc_6_input_sync_blk[3] | proc_6_output_sync_blk[3]);
    assign proc_6_data_FIFO_blk[4] = 1'b0;
    assign proc_6_data_PIPO_blk[4] = 1'b0;
    assign proc_6_start_FIFO_blk[4] = 1'b0;
    assign proc_6_TLF_FIFO_blk[4] = 1'b0;
    assign proc_6_input_sync_blk[4] = 1'b0 | (ap_sync_load_value35_U0_ap_ready & load_value35_U0.ap_idle & ~ap_sync_load_value32_U0_ap_ready);
    assign proc_6_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_6[4] = dl_detect_out ? proc_dep_vld_vec_6_reg[4] : (proc_6_data_FIFO_blk[4] | proc_6_data_PIPO_blk[4] | proc_6_start_FIFO_blk[4] | proc_6_TLF_FIFO_blk[4] | proc_6_input_sync_blk[4] | proc_6_output_sync_blk[4]);
    assign proc_6_data_FIFO_blk[5] = 1'b0;
    assign proc_6_data_PIPO_blk[5] = 1'b0;
    assign proc_6_start_FIFO_blk[5] = 1'b0;
    assign proc_6_TLF_FIFO_blk[5] = 1'b0;
    assign proc_6_input_sync_blk[5] = 1'b0 | (ap_sync_load_value35_U0_ap_ready & load_value35_U0.ap_idle & ~ap_sync_load_value33_U0_ap_ready);
    assign proc_6_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_6[5] = dl_detect_out ? proc_dep_vld_vec_6_reg[5] : (proc_6_data_FIFO_blk[5] | proc_6_data_PIPO_blk[5] | proc_6_start_FIFO_blk[5] | proc_6_TLF_FIFO_blk[5] | proc_6_input_sync_blk[5] | proc_6_output_sync_blk[5]);
    assign proc_6_data_FIFO_blk[6] = 1'b0;
    assign proc_6_data_PIPO_blk[6] = 1'b0;
    assign proc_6_start_FIFO_blk[6] = 1'b0;
    assign proc_6_TLF_FIFO_blk[6] = 1'b0;
    assign proc_6_input_sync_blk[6] = 1'b0 | (ap_sync_load_value35_U0_ap_ready & load_value35_U0.ap_idle & ~ap_sync_load_value34_U0_ap_ready);
    assign proc_6_output_sync_blk[6] = 1'b0;
    assign proc_dep_vld_vec_6[6] = dl_detect_out ? proc_dep_vld_vec_6_reg[6] : (proc_6_data_FIFO_blk[6] | proc_6_data_PIPO_blk[6] | proc_6_start_FIFO_blk[6] | proc_6_TLF_FIFO_blk[6] | proc_6_input_sync_blk[6] | proc_6_output_sync_blk[6]);
    assign proc_6_data_FIFO_blk[7] = 1'b0;
    assign proc_6_data_PIPO_blk[7] = 1'b0;
    assign proc_6_start_FIFO_blk[7] = 1'b0;
    assign proc_6_TLF_FIFO_blk[7] = 1'b0;
    assign proc_6_input_sync_blk[7] = 1'b0 | (ap_sync_load_value35_U0_ap_ready & load_value35_U0.ap_idle & ~ap_sync_load_value36_U0_ap_ready);
    assign proc_6_output_sync_blk[7] = 1'b0;
    assign proc_dep_vld_vec_6[7] = dl_detect_out ? proc_dep_vld_vec_6_reg[7] : (proc_6_data_FIFO_blk[7] | proc_6_data_PIPO_blk[7] | proc_6_start_FIFO_blk[7] | proc_6_TLF_FIFO_blk[7] | proc_6_input_sync_blk[7] | proc_6_output_sync_blk[7]);
    assign proc_6_data_FIFO_blk[8] = 1'b0;
    assign proc_6_data_PIPO_blk[8] = 1'b0;
    assign proc_6_start_FIFO_blk[8] = 1'b0;
    assign proc_6_TLF_FIFO_blk[8] = 1'b0;
    assign proc_6_input_sync_blk[8] = 1'b0 | (ap_sync_load_value35_U0_ap_ready & load_value35_U0.ap_idle & ~ap_sync_load_value37_U0_ap_ready);
    assign proc_6_output_sync_blk[8] = 1'b0;
    assign proc_dep_vld_vec_6[8] = dl_detect_out ? proc_dep_vld_vec_6_reg[8] : (proc_6_data_FIFO_blk[8] | proc_6_data_PIPO_blk[8] | proc_6_start_FIFO_blk[8] | proc_6_TLF_FIFO_blk[8] | proc_6_input_sync_blk[8] | proc_6_output_sync_blk[8]);
    assign proc_6_data_FIFO_blk[9] = 1'b0;
    assign proc_6_data_PIPO_blk[9] = 1'b0;
    assign proc_6_start_FIFO_blk[9] = 1'b0;
    assign proc_6_TLF_FIFO_blk[9] = 1'b0;
    assign proc_6_input_sync_blk[9] = 1'b0 | (ap_sync_load_value35_U0_ap_ready & load_value35_U0.ap_idle & ~ap_sync_load_value38_U0_ap_ready);
    assign proc_6_output_sync_blk[9] = 1'b0;
    assign proc_dep_vld_vec_6[9] = dl_detect_out ? proc_dep_vld_vec_6_reg[9] : (proc_6_data_FIFO_blk[9] | proc_6_data_PIPO_blk[9] | proc_6_start_FIFO_blk[9] | proc_6_TLF_FIFO_blk[9] | proc_6_input_sync_blk[9] | proc_6_output_sync_blk[9]);
    assign proc_6_data_FIFO_blk[10] = 1'b0;
    assign proc_6_data_PIPO_blk[10] = 1'b0;
    assign proc_6_start_FIFO_blk[10] = 1'b0;
    assign proc_6_TLF_FIFO_blk[10] = 1'b0;
    assign proc_6_input_sync_blk[10] = 1'b0 | (ap_sync_load_value35_U0_ap_ready & load_value35_U0.ap_idle & ~ap_sync_load_value39_U0_ap_ready);
    assign proc_6_output_sync_blk[10] = 1'b0;
    assign proc_dep_vld_vec_6[10] = dl_detect_out ? proc_dep_vld_vec_6_reg[10] : (proc_6_data_FIFO_blk[10] | proc_6_data_PIPO_blk[10] | proc_6_start_FIFO_blk[10] | proc_6_TLF_FIFO_blk[10] | proc_6_input_sync_blk[10] | proc_6_output_sync_blk[10]);
    assign proc_6_data_FIFO_blk[11] = 1'b0;
    assign proc_6_data_PIPO_blk[11] = 1'b0;
    assign proc_6_start_FIFO_blk[11] = 1'b0;
    assign proc_6_TLF_FIFO_blk[11] = 1'b0;
    assign proc_6_input_sync_blk[11] = 1'b0 | (ap_sync_load_value35_U0_ap_ready & load_value35_U0.ap_idle & ~ap_sync_load_value40_U0_ap_ready);
    assign proc_6_output_sync_blk[11] = 1'b0;
    assign proc_dep_vld_vec_6[11] = dl_detect_out ? proc_dep_vld_vec_6_reg[11] : (proc_6_data_FIFO_blk[11] | proc_6_data_PIPO_blk[11] | proc_6_start_FIFO_blk[11] | proc_6_TLF_FIFO_blk[11] | proc_6_input_sync_blk[11] | proc_6_output_sync_blk[11]);
    assign proc_6_data_FIFO_blk[12] = 1'b0;
    assign proc_6_data_PIPO_blk[12] = 1'b0;
    assign proc_6_start_FIFO_blk[12] = 1'b0;
    assign proc_6_TLF_FIFO_blk[12] = 1'b0;
    assign proc_6_input_sync_blk[12] = 1'b0 | (ap_sync_load_value35_U0_ap_ready & load_value35_U0.ap_idle & ~ap_sync_load_value41_U0_ap_ready);
    assign proc_6_output_sync_blk[12] = 1'b0;
    assign proc_dep_vld_vec_6[12] = dl_detect_out ? proc_dep_vld_vec_6_reg[12] : (proc_6_data_FIFO_blk[12] | proc_6_data_PIPO_blk[12] | proc_6_start_FIFO_blk[12] | proc_6_TLF_FIFO_blk[12] | proc_6_input_sync_blk[12] | proc_6_output_sync_blk[12]);
    assign proc_6_data_FIFO_blk[13] = 1'b0;
    assign proc_6_data_PIPO_blk[13] = 1'b0;
    assign proc_6_start_FIFO_blk[13] = 1'b0;
    assign proc_6_TLF_FIFO_blk[13] = 1'b0;
    assign proc_6_input_sync_blk[13] = 1'b0 | (ap_sync_load_value35_U0_ap_ready & load_value35_U0.ap_idle & ~ap_sync_load_value42_U0_ap_ready);
    assign proc_6_output_sync_blk[13] = 1'b0;
    assign proc_dep_vld_vec_6[13] = dl_detect_out ? proc_dep_vld_vec_6_reg[13] : (proc_6_data_FIFO_blk[13] | proc_6_data_PIPO_blk[13] | proc_6_start_FIFO_blk[13] | proc_6_TLF_FIFO_blk[13] | proc_6_input_sync_blk[13] | proc_6_output_sync_blk[13]);
    assign proc_6_data_FIFO_blk[14] = 1'b0;
    assign proc_6_data_PIPO_blk[14] = 1'b0;
    assign proc_6_start_FIFO_blk[14] = 1'b0;
    assign proc_6_TLF_FIFO_blk[14] = 1'b0;
    assign proc_6_input_sync_blk[14] = 1'b0 | (ap_sync_load_value35_U0_ap_ready & load_value35_U0.ap_idle & ~ap_sync_load_value43_U0_ap_ready);
    assign proc_6_output_sync_blk[14] = 1'b0;
    assign proc_dep_vld_vec_6[14] = dl_detect_out ? proc_dep_vld_vec_6_reg[14] : (proc_6_data_FIFO_blk[14] | proc_6_data_PIPO_blk[14] | proc_6_start_FIFO_blk[14] | proc_6_TLF_FIFO_blk[14] | proc_6_input_sync_blk[14] | proc_6_output_sync_blk[14]);
    assign proc_6_data_FIFO_blk[15] = 1'b0;
    assign proc_6_data_PIPO_blk[15] = 1'b0;
    assign proc_6_start_FIFO_blk[15] = 1'b0;
    assign proc_6_TLF_FIFO_blk[15] = 1'b0;
    assign proc_6_input_sync_blk[15] = 1'b0 | (ap_sync_load_value35_U0_ap_ready & load_value35_U0.ap_idle & ~ap_sync_load_value44_U0_ap_ready);
    assign proc_6_output_sync_blk[15] = 1'b0;
    assign proc_dep_vld_vec_6[15] = dl_detect_out ? proc_dep_vld_vec_6_reg[15] : (proc_6_data_FIFO_blk[15] | proc_6_data_PIPO_blk[15] | proc_6_start_FIFO_blk[15] | proc_6_TLF_FIFO_blk[15] | proc_6_input_sync_blk[15] | proc_6_output_sync_blk[15]);
    assign proc_6_data_FIFO_blk[16] = 1'b0;
    assign proc_6_data_PIPO_blk[16] = 1'b0;
    assign proc_6_start_FIFO_blk[16] = 1'b0;
    assign proc_6_TLF_FIFO_blk[16] = 1'b0;
    assign proc_6_input_sync_blk[16] = 1'b0 | (ap_sync_load_value35_U0_ap_ready & load_value35_U0.ap_idle & ~ap_sync_load_value45_U0_ap_ready);
    assign proc_6_output_sync_blk[16] = 1'b0;
    assign proc_dep_vld_vec_6[16] = dl_detect_out ? proc_dep_vld_vec_6_reg[16] : (proc_6_data_FIFO_blk[16] | proc_6_data_PIPO_blk[16] | proc_6_start_FIFO_blk[16] | proc_6_TLF_FIFO_blk[16] | proc_6_input_sync_blk[16] | proc_6_output_sync_blk[16]);
    assign proc_6_data_FIFO_blk[17] = 1'b0;
    assign proc_6_data_PIPO_blk[17] = 1'b0;
    assign proc_6_start_FIFO_blk[17] = 1'b0;
    assign proc_6_TLF_FIFO_blk[17] = 1'b0;
    assign proc_6_input_sync_blk[17] = 1'b0 | (ap_sync_load_value35_U0_ap_ready & load_value35_U0.ap_idle & ~ap_sync_load_value46_U0_ap_ready);
    assign proc_6_output_sync_blk[17] = 1'b0;
    assign proc_dep_vld_vec_6[17] = dl_detect_out ? proc_dep_vld_vec_6_reg[17] : (proc_6_data_FIFO_blk[17] | proc_6_data_PIPO_blk[17] | proc_6_start_FIFO_blk[17] | proc_6_TLF_FIFO_blk[17] | proc_6_input_sync_blk[17] | proc_6_output_sync_blk[17]);
    assign proc_6_data_FIFO_blk[18] = 1'b0;
    assign proc_6_data_PIPO_blk[18] = 1'b0;
    assign proc_6_start_FIFO_blk[18] = 1'b0;
    assign proc_6_TLF_FIFO_blk[18] = 1'b0;
    assign proc_6_input_sync_blk[18] = 1'b0 | (ap_sync_load_value35_U0_ap_ready & load_value35_U0.ap_idle & ~ap_sync_load_value47_U0_ap_ready);
    assign proc_6_output_sync_blk[18] = 1'b0;
    assign proc_dep_vld_vec_6[18] = dl_detect_out ? proc_dep_vld_vec_6_reg[18] : (proc_6_data_FIFO_blk[18] | proc_6_data_PIPO_blk[18] | proc_6_start_FIFO_blk[18] | proc_6_TLF_FIFO_blk[18] | proc_6_input_sync_blk[18] | proc_6_output_sync_blk[18]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_6_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_6_reg <= proc_dep_vld_vec_6;
        end
    end
    assign in_chan_dep_vld_vec_6[0] = dep_chan_vld_0_6;
    assign in_chan_dep_data_vec_6[34 : 0] = dep_chan_data_0_6;
    assign token_in_vec_6[0] = token_0_6;
    assign in_chan_dep_vld_vec_6[1] = dep_chan_vld_1_6;
    assign in_chan_dep_data_vec_6[69 : 35] = dep_chan_data_1_6;
    assign token_in_vec_6[1] = token_1_6;
    assign in_chan_dep_vld_vec_6[2] = dep_chan_vld_2_6;
    assign in_chan_dep_data_vec_6[104 : 70] = dep_chan_data_2_6;
    assign token_in_vec_6[2] = token_2_6;
    assign in_chan_dep_vld_vec_6[3] = dep_chan_vld_3_6;
    assign in_chan_dep_data_vec_6[139 : 105] = dep_chan_data_3_6;
    assign token_in_vec_6[3] = token_3_6;
    assign in_chan_dep_vld_vec_6[4] = dep_chan_vld_4_6;
    assign in_chan_dep_data_vec_6[174 : 140] = dep_chan_data_4_6;
    assign token_in_vec_6[4] = token_4_6;
    assign in_chan_dep_vld_vec_6[5] = dep_chan_vld_5_6;
    assign in_chan_dep_data_vec_6[209 : 175] = dep_chan_data_5_6;
    assign token_in_vec_6[5] = token_5_6;
    assign in_chan_dep_vld_vec_6[6] = dep_chan_vld_7_6;
    assign in_chan_dep_data_vec_6[244 : 210] = dep_chan_data_7_6;
    assign token_in_vec_6[6] = token_7_6;
    assign in_chan_dep_vld_vec_6[7] = dep_chan_vld_8_6;
    assign in_chan_dep_data_vec_6[279 : 245] = dep_chan_data_8_6;
    assign token_in_vec_6[7] = token_8_6;
    assign in_chan_dep_vld_vec_6[8] = dep_chan_vld_9_6;
    assign in_chan_dep_data_vec_6[314 : 280] = dep_chan_data_9_6;
    assign token_in_vec_6[8] = token_9_6;
    assign in_chan_dep_vld_vec_6[9] = dep_chan_vld_10_6;
    assign in_chan_dep_data_vec_6[349 : 315] = dep_chan_data_10_6;
    assign token_in_vec_6[9] = token_10_6;
    assign in_chan_dep_vld_vec_6[10] = dep_chan_vld_11_6;
    assign in_chan_dep_data_vec_6[384 : 350] = dep_chan_data_11_6;
    assign token_in_vec_6[10] = token_11_6;
    assign in_chan_dep_vld_vec_6[11] = dep_chan_vld_12_6;
    assign in_chan_dep_data_vec_6[419 : 385] = dep_chan_data_12_6;
    assign token_in_vec_6[11] = token_12_6;
    assign in_chan_dep_vld_vec_6[12] = dep_chan_vld_13_6;
    assign in_chan_dep_data_vec_6[454 : 420] = dep_chan_data_13_6;
    assign token_in_vec_6[12] = token_13_6;
    assign in_chan_dep_vld_vec_6[13] = dep_chan_vld_14_6;
    assign in_chan_dep_data_vec_6[489 : 455] = dep_chan_data_14_6;
    assign token_in_vec_6[13] = token_14_6;
    assign in_chan_dep_vld_vec_6[14] = dep_chan_vld_15_6;
    assign in_chan_dep_data_vec_6[524 : 490] = dep_chan_data_15_6;
    assign token_in_vec_6[14] = token_15_6;
    assign in_chan_dep_vld_vec_6[15] = dep_chan_vld_16_6;
    assign in_chan_dep_data_vec_6[559 : 525] = dep_chan_data_16_6;
    assign token_in_vec_6[15] = token_16_6;
    assign in_chan_dep_vld_vec_6[16] = dep_chan_vld_17_6;
    assign in_chan_dep_data_vec_6[594 : 560] = dep_chan_data_17_6;
    assign token_in_vec_6[16] = token_17_6;
    assign in_chan_dep_vld_vec_6[17] = dep_chan_vld_18_6;
    assign in_chan_dep_data_vec_6[629 : 595] = dep_chan_data_18_6;
    assign token_in_vec_6[17] = token_18_6;
    assign in_chan_dep_vld_vec_6[18] = dep_chan_vld_22_6;
    assign in_chan_dep_data_vec_6[664 : 630] = dep_chan_data_22_6;
    assign token_in_vec_6[18] = token_22_6;
    assign dep_chan_vld_6_0 = out_chan_dep_vld_vec_6[0];
    assign dep_chan_data_6_0 = out_chan_dep_data_6;
    assign token_6_0 = token_out_vec_6[0];
    assign dep_chan_vld_6_1 = out_chan_dep_vld_vec_6[1];
    assign dep_chan_data_6_1 = out_chan_dep_data_6;
    assign token_6_1 = token_out_vec_6[1];
    assign dep_chan_vld_6_22 = out_chan_dep_vld_vec_6[2];
    assign dep_chan_data_6_22 = out_chan_dep_data_6;
    assign token_6_22 = token_out_vec_6[2];
    assign dep_chan_vld_6_2 = out_chan_dep_vld_vec_6[3];
    assign dep_chan_data_6_2 = out_chan_dep_data_6;
    assign token_6_2 = token_out_vec_6[3];
    assign dep_chan_vld_6_3 = out_chan_dep_vld_vec_6[4];
    assign dep_chan_data_6_3 = out_chan_dep_data_6;
    assign token_6_3 = token_out_vec_6[4];
    assign dep_chan_vld_6_4 = out_chan_dep_vld_vec_6[5];
    assign dep_chan_data_6_4 = out_chan_dep_data_6;
    assign token_6_4 = token_out_vec_6[5];
    assign dep_chan_vld_6_5 = out_chan_dep_vld_vec_6[6];
    assign dep_chan_data_6_5 = out_chan_dep_data_6;
    assign token_6_5 = token_out_vec_6[6];
    assign dep_chan_vld_6_7 = out_chan_dep_vld_vec_6[7];
    assign dep_chan_data_6_7 = out_chan_dep_data_6;
    assign token_6_7 = token_out_vec_6[7];
    assign dep_chan_vld_6_8 = out_chan_dep_vld_vec_6[8];
    assign dep_chan_data_6_8 = out_chan_dep_data_6;
    assign token_6_8 = token_out_vec_6[8];
    assign dep_chan_vld_6_9 = out_chan_dep_vld_vec_6[9];
    assign dep_chan_data_6_9 = out_chan_dep_data_6;
    assign token_6_9 = token_out_vec_6[9];
    assign dep_chan_vld_6_10 = out_chan_dep_vld_vec_6[10];
    assign dep_chan_data_6_10 = out_chan_dep_data_6;
    assign token_6_10 = token_out_vec_6[10];
    assign dep_chan_vld_6_11 = out_chan_dep_vld_vec_6[11];
    assign dep_chan_data_6_11 = out_chan_dep_data_6;
    assign token_6_11 = token_out_vec_6[11];
    assign dep_chan_vld_6_12 = out_chan_dep_vld_vec_6[12];
    assign dep_chan_data_6_12 = out_chan_dep_data_6;
    assign token_6_12 = token_out_vec_6[12];
    assign dep_chan_vld_6_13 = out_chan_dep_vld_vec_6[13];
    assign dep_chan_data_6_13 = out_chan_dep_data_6;
    assign token_6_13 = token_out_vec_6[13];
    assign dep_chan_vld_6_14 = out_chan_dep_vld_vec_6[14];
    assign dep_chan_data_6_14 = out_chan_dep_data_6;
    assign token_6_14 = token_out_vec_6[14];
    assign dep_chan_vld_6_15 = out_chan_dep_vld_vec_6[15];
    assign dep_chan_data_6_15 = out_chan_dep_data_6;
    assign token_6_15 = token_out_vec_6[15];
    assign dep_chan_vld_6_16 = out_chan_dep_vld_vec_6[16];
    assign dep_chan_data_6_16 = out_chan_dep_data_6;
    assign token_6_16 = token_out_vec_6[16];
    assign dep_chan_vld_6_17 = out_chan_dep_vld_vec_6[17];
    assign dep_chan_data_6_17 = out_chan_dep_data_6;
    assign token_6_17 = token_out_vec_6[17];
    assign dep_chan_vld_6_18 = out_chan_dep_vld_vec_6[18];
    assign dep_chan_data_6_18 = out_chan_dep_data_6;
    assign token_6_18 = token_out_vec_6[18];

    // Process: load_value36_U0
    kernel_pr_hls_deadlock_detect_unit #(35, 7, 19, 19) kernel_pr_hls_deadlock_detect_unit_7 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_7),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_7),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_7),
        .token_in_vec(token_in_vec_7),
        .dl_detect_in(dl_detect_out),
        .origin(origin[7]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_7),
        .out_chan_dep_data(out_chan_dep_data_7),
        .token_out_vec(token_out_vec_7),
        .dl_detect_out(dl_in_vec[7]));

    assign proc_7_data_FIFO_blk[0] = 1'b0 | (~load_value36_U0.value_r_blk_n);
    assign proc_7_data_PIPO_blk[0] = 1'b0;
    assign proc_7_start_FIFO_blk[0] = 1'b0;
    assign proc_7_TLF_FIFO_blk[0] = 1'b0;
    assign proc_7_input_sync_blk[0] = 1'b0 | (ap_sync_load_value36_U0_ap_ready & load_value36_U0.ap_idle & ~ap_sync_kernel_pr_entry98_U0_ap_ready);
    assign proc_7_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_7[0] = dl_detect_out ? proc_dep_vld_vec_7_reg[0] : (proc_7_data_FIFO_blk[0] | proc_7_data_PIPO_blk[0] | proc_7_start_FIFO_blk[0] | proc_7_TLF_FIFO_blk[0] | proc_7_input_sync_blk[0] | proc_7_output_sync_blk[0]);
    assign proc_7_data_FIFO_blk[1] = 1'b0 | (~load_value36_U0.bipedge_size_blk_n) | (~load_value36_U0.bipedge_stream_V_V4_blk_n);
    assign proc_7_data_PIPO_blk[1] = 1'b0;
    assign proc_7_start_FIFO_blk[1] = 1'b0;
    assign proc_7_TLF_FIFO_blk[1] = 1'b0;
    assign proc_7_input_sync_blk[1] = 1'b0 | (ap_sync_load_value36_U0_ap_ready & load_value36_U0.ap_idle & ~ap_sync_load_bipedge30_U0_ap_ready);
    assign proc_7_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_7[1] = dl_detect_out ? proc_dep_vld_vec_7_reg[1] : (proc_7_data_FIFO_blk[1] | proc_7_data_PIPO_blk[1] | proc_7_start_FIFO_blk[1] | proc_7_TLF_FIFO_blk[1] | proc_7_input_sync_blk[1] | proc_7_output_sync_blk[1]);
    assign proc_7_data_FIFO_blk[2] = 1'b0 | (~load_value36_U0.value_stream_V_V19_blk_n);
    assign proc_7_data_PIPO_blk[2] = 1'b0;
    assign proc_7_start_FIFO_blk[2] = 1'b0;
    assign proc_7_TLF_FIFO_blk[2] = 1'b0;
    assign proc_7_input_sync_blk[2] = 1'b0;
    assign proc_7_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_7[2] = dl_detect_out ? proc_dep_vld_vec_7_reg[2] : (proc_7_data_FIFO_blk[2] | proc_7_data_PIPO_blk[2] | proc_7_start_FIFO_blk[2] | proc_7_TLF_FIFO_blk[2] | proc_7_input_sync_blk[2] | proc_7_output_sync_blk[2]);
    assign proc_7_data_FIFO_blk[3] = 1'b0;
    assign proc_7_data_PIPO_blk[3] = 1'b0;
    assign proc_7_start_FIFO_blk[3] = 1'b0;
    assign proc_7_TLF_FIFO_blk[3] = 1'b0;
    assign proc_7_input_sync_blk[3] = 1'b0 | (ap_sync_load_value36_U0_ap_ready & load_value36_U0.ap_idle & ~ap_sync_load_bipedge31_U0_ap_ready);
    assign proc_7_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_7[3] = dl_detect_out ? proc_dep_vld_vec_7_reg[3] : (proc_7_data_FIFO_blk[3] | proc_7_data_PIPO_blk[3] | proc_7_start_FIFO_blk[3] | proc_7_TLF_FIFO_blk[3] | proc_7_input_sync_blk[3] | proc_7_output_sync_blk[3]);
    assign proc_7_data_FIFO_blk[4] = 1'b0;
    assign proc_7_data_PIPO_blk[4] = 1'b0;
    assign proc_7_start_FIFO_blk[4] = 1'b0;
    assign proc_7_TLF_FIFO_blk[4] = 1'b0;
    assign proc_7_input_sync_blk[4] = 1'b0 | (ap_sync_load_value36_U0_ap_ready & load_value36_U0.ap_idle & ~ap_sync_load_value32_U0_ap_ready);
    assign proc_7_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_7[4] = dl_detect_out ? proc_dep_vld_vec_7_reg[4] : (proc_7_data_FIFO_blk[4] | proc_7_data_PIPO_blk[4] | proc_7_start_FIFO_blk[4] | proc_7_TLF_FIFO_blk[4] | proc_7_input_sync_blk[4] | proc_7_output_sync_blk[4]);
    assign proc_7_data_FIFO_blk[5] = 1'b0;
    assign proc_7_data_PIPO_blk[5] = 1'b0;
    assign proc_7_start_FIFO_blk[5] = 1'b0;
    assign proc_7_TLF_FIFO_blk[5] = 1'b0;
    assign proc_7_input_sync_blk[5] = 1'b0 | (ap_sync_load_value36_U0_ap_ready & load_value36_U0.ap_idle & ~ap_sync_load_value33_U0_ap_ready);
    assign proc_7_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_7[5] = dl_detect_out ? proc_dep_vld_vec_7_reg[5] : (proc_7_data_FIFO_blk[5] | proc_7_data_PIPO_blk[5] | proc_7_start_FIFO_blk[5] | proc_7_TLF_FIFO_blk[5] | proc_7_input_sync_blk[5] | proc_7_output_sync_blk[5]);
    assign proc_7_data_FIFO_blk[6] = 1'b0;
    assign proc_7_data_PIPO_blk[6] = 1'b0;
    assign proc_7_start_FIFO_blk[6] = 1'b0;
    assign proc_7_TLF_FIFO_blk[6] = 1'b0;
    assign proc_7_input_sync_blk[6] = 1'b0 | (ap_sync_load_value36_U0_ap_ready & load_value36_U0.ap_idle & ~ap_sync_load_value34_U0_ap_ready);
    assign proc_7_output_sync_blk[6] = 1'b0;
    assign proc_dep_vld_vec_7[6] = dl_detect_out ? proc_dep_vld_vec_7_reg[6] : (proc_7_data_FIFO_blk[6] | proc_7_data_PIPO_blk[6] | proc_7_start_FIFO_blk[6] | proc_7_TLF_FIFO_blk[6] | proc_7_input_sync_blk[6] | proc_7_output_sync_blk[6]);
    assign proc_7_data_FIFO_blk[7] = 1'b0;
    assign proc_7_data_PIPO_blk[7] = 1'b0;
    assign proc_7_start_FIFO_blk[7] = 1'b0;
    assign proc_7_TLF_FIFO_blk[7] = 1'b0;
    assign proc_7_input_sync_blk[7] = 1'b0 | (ap_sync_load_value36_U0_ap_ready & load_value36_U0.ap_idle & ~ap_sync_load_value35_U0_ap_ready);
    assign proc_7_output_sync_blk[7] = 1'b0;
    assign proc_dep_vld_vec_7[7] = dl_detect_out ? proc_dep_vld_vec_7_reg[7] : (proc_7_data_FIFO_blk[7] | proc_7_data_PIPO_blk[7] | proc_7_start_FIFO_blk[7] | proc_7_TLF_FIFO_blk[7] | proc_7_input_sync_blk[7] | proc_7_output_sync_blk[7]);
    assign proc_7_data_FIFO_blk[8] = 1'b0;
    assign proc_7_data_PIPO_blk[8] = 1'b0;
    assign proc_7_start_FIFO_blk[8] = 1'b0;
    assign proc_7_TLF_FIFO_blk[8] = 1'b0;
    assign proc_7_input_sync_blk[8] = 1'b0 | (ap_sync_load_value36_U0_ap_ready & load_value36_U0.ap_idle & ~ap_sync_load_value37_U0_ap_ready);
    assign proc_7_output_sync_blk[8] = 1'b0;
    assign proc_dep_vld_vec_7[8] = dl_detect_out ? proc_dep_vld_vec_7_reg[8] : (proc_7_data_FIFO_blk[8] | proc_7_data_PIPO_blk[8] | proc_7_start_FIFO_blk[8] | proc_7_TLF_FIFO_blk[8] | proc_7_input_sync_blk[8] | proc_7_output_sync_blk[8]);
    assign proc_7_data_FIFO_blk[9] = 1'b0;
    assign proc_7_data_PIPO_blk[9] = 1'b0;
    assign proc_7_start_FIFO_blk[9] = 1'b0;
    assign proc_7_TLF_FIFO_blk[9] = 1'b0;
    assign proc_7_input_sync_blk[9] = 1'b0 | (ap_sync_load_value36_U0_ap_ready & load_value36_U0.ap_idle & ~ap_sync_load_value38_U0_ap_ready);
    assign proc_7_output_sync_blk[9] = 1'b0;
    assign proc_dep_vld_vec_7[9] = dl_detect_out ? proc_dep_vld_vec_7_reg[9] : (proc_7_data_FIFO_blk[9] | proc_7_data_PIPO_blk[9] | proc_7_start_FIFO_blk[9] | proc_7_TLF_FIFO_blk[9] | proc_7_input_sync_blk[9] | proc_7_output_sync_blk[9]);
    assign proc_7_data_FIFO_blk[10] = 1'b0;
    assign proc_7_data_PIPO_blk[10] = 1'b0;
    assign proc_7_start_FIFO_blk[10] = 1'b0;
    assign proc_7_TLF_FIFO_blk[10] = 1'b0;
    assign proc_7_input_sync_blk[10] = 1'b0 | (ap_sync_load_value36_U0_ap_ready & load_value36_U0.ap_idle & ~ap_sync_load_value39_U0_ap_ready);
    assign proc_7_output_sync_blk[10] = 1'b0;
    assign proc_dep_vld_vec_7[10] = dl_detect_out ? proc_dep_vld_vec_7_reg[10] : (proc_7_data_FIFO_blk[10] | proc_7_data_PIPO_blk[10] | proc_7_start_FIFO_blk[10] | proc_7_TLF_FIFO_blk[10] | proc_7_input_sync_blk[10] | proc_7_output_sync_blk[10]);
    assign proc_7_data_FIFO_blk[11] = 1'b0;
    assign proc_7_data_PIPO_blk[11] = 1'b0;
    assign proc_7_start_FIFO_blk[11] = 1'b0;
    assign proc_7_TLF_FIFO_blk[11] = 1'b0;
    assign proc_7_input_sync_blk[11] = 1'b0 | (ap_sync_load_value36_U0_ap_ready & load_value36_U0.ap_idle & ~ap_sync_load_value40_U0_ap_ready);
    assign proc_7_output_sync_blk[11] = 1'b0;
    assign proc_dep_vld_vec_7[11] = dl_detect_out ? proc_dep_vld_vec_7_reg[11] : (proc_7_data_FIFO_blk[11] | proc_7_data_PIPO_blk[11] | proc_7_start_FIFO_blk[11] | proc_7_TLF_FIFO_blk[11] | proc_7_input_sync_blk[11] | proc_7_output_sync_blk[11]);
    assign proc_7_data_FIFO_blk[12] = 1'b0;
    assign proc_7_data_PIPO_blk[12] = 1'b0;
    assign proc_7_start_FIFO_blk[12] = 1'b0;
    assign proc_7_TLF_FIFO_blk[12] = 1'b0;
    assign proc_7_input_sync_blk[12] = 1'b0 | (ap_sync_load_value36_U0_ap_ready & load_value36_U0.ap_idle & ~ap_sync_load_value41_U0_ap_ready);
    assign proc_7_output_sync_blk[12] = 1'b0;
    assign proc_dep_vld_vec_7[12] = dl_detect_out ? proc_dep_vld_vec_7_reg[12] : (proc_7_data_FIFO_blk[12] | proc_7_data_PIPO_blk[12] | proc_7_start_FIFO_blk[12] | proc_7_TLF_FIFO_blk[12] | proc_7_input_sync_blk[12] | proc_7_output_sync_blk[12]);
    assign proc_7_data_FIFO_blk[13] = 1'b0;
    assign proc_7_data_PIPO_blk[13] = 1'b0;
    assign proc_7_start_FIFO_blk[13] = 1'b0;
    assign proc_7_TLF_FIFO_blk[13] = 1'b0;
    assign proc_7_input_sync_blk[13] = 1'b0 | (ap_sync_load_value36_U0_ap_ready & load_value36_U0.ap_idle & ~ap_sync_load_value42_U0_ap_ready);
    assign proc_7_output_sync_blk[13] = 1'b0;
    assign proc_dep_vld_vec_7[13] = dl_detect_out ? proc_dep_vld_vec_7_reg[13] : (proc_7_data_FIFO_blk[13] | proc_7_data_PIPO_blk[13] | proc_7_start_FIFO_blk[13] | proc_7_TLF_FIFO_blk[13] | proc_7_input_sync_blk[13] | proc_7_output_sync_blk[13]);
    assign proc_7_data_FIFO_blk[14] = 1'b0;
    assign proc_7_data_PIPO_blk[14] = 1'b0;
    assign proc_7_start_FIFO_blk[14] = 1'b0;
    assign proc_7_TLF_FIFO_blk[14] = 1'b0;
    assign proc_7_input_sync_blk[14] = 1'b0 | (ap_sync_load_value36_U0_ap_ready & load_value36_U0.ap_idle & ~ap_sync_load_value43_U0_ap_ready);
    assign proc_7_output_sync_blk[14] = 1'b0;
    assign proc_dep_vld_vec_7[14] = dl_detect_out ? proc_dep_vld_vec_7_reg[14] : (proc_7_data_FIFO_blk[14] | proc_7_data_PIPO_blk[14] | proc_7_start_FIFO_blk[14] | proc_7_TLF_FIFO_blk[14] | proc_7_input_sync_blk[14] | proc_7_output_sync_blk[14]);
    assign proc_7_data_FIFO_blk[15] = 1'b0;
    assign proc_7_data_PIPO_blk[15] = 1'b0;
    assign proc_7_start_FIFO_blk[15] = 1'b0;
    assign proc_7_TLF_FIFO_blk[15] = 1'b0;
    assign proc_7_input_sync_blk[15] = 1'b0 | (ap_sync_load_value36_U0_ap_ready & load_value36_U0.ap_idle & ~ap_sync_load_value44_U0_ap_ready);
    assign proc_7_output_sync_blk[15] = 1'b0;
    assign proc_dep_vld_vec_7[15] = dl_detect_out ? proc_dep_vld_vec_7_reg[15] : (proc_7_data_FIFO_blk[15] | proc_7_data_PIPO_blk[15] | proc_7_start_FIFO_blk[15] | proc_7_TLF_FIFO_blk[15] | proc_7_input_sync_blk[15] | proc_7_output_sync_blk[15]);
    assign proc_7_data_FIFO_blk[16] = 1'b0;
    assign proc_7_data_PIPO_blk[16] = 1'b0;
    assign proc_7_start_FIFO_blk[16] = 1'b0;
    assign proc_7_TLF_FIFO_blk[16] = 1'b0;
    assign proc_7_input_sync_blk[16] = 1'b0 | (ap_sync_load_value36_U0_ap_ready & load_value36_U0.ap_idle & ~ap_sync_load_value45_U0_ap_ready);
    assign proc_7_output_sync_blk[16] = 1'b0;
    assign proc_dep_vld_vec_7[16] = dl_detect_out ? proc_dep_vld_vec_7_reg[16] : (proc_7_data_FIFO_blk[16] | proc_7_data_PIPO_blk[16] | proc_7_start_FIFO_blk[16] | proc_7_TLF_FIFO_blk[16] | proc_7_input_sync_blk[16] | proc_7_output_sync_blk[16]);
    assign proc_7_data_FIFO_blk[17] = 1'b0;
    assign proc_7_data_PIPO_blk[17] = 1'b0;
    assign proc_7_start_FIFO_blk[17] = 1'b0;
    assign proc_7_TLF_FIFO_blk[17] = 1'b0;
    assign proc_7_input_sync_blk[17] = 1'b0 | (ap_sync_load_value36_U0_ap_ready & load_value36_U0.ap_idle & ~ap_sync_load_value46_U0_ap_ready);
    assign proc_7_output_sync_blk[17] = 1'b0;
    assign proc_dep_vld_vec_7[17] = dl_detect_out ? proc_dep_vld_vec_7_reg[17] : (proc_7_data_FIFO_blk[17] | proc_7_data_PIPO_blk[17] | proc_7_start_FIFO_blk[17] | proc_7_TLF_FIFO_blk[17] | proc_7_input_sync_blk[17] | proc_7_output_sync_blk[17]);
    assign proc_7_data_FIFO_blk[18] = 1'b0;
    assign proc_7_data_PIPO_blk[18] = 1'b0;
    assign proc_7_start_FIFO_blk[18] = 1'b0;
    assign proc_7_TLF_FIFO_blk[18] = 1'b0;
    assign proc_7_input_sync_blk[18] = 1'b0 | (ap_sync_load_value36_U0_ap_ready & load_value36_U0.ap_idle & ~ap_sync_load_value47_U0_ap_ready);
    assign proc_7_output_sync_blk[18] = 1'b0;
    assign proc_dep_vld_vec_7[18] = dl_detect_out ? proc_dep_vld_vec_7_reg[18] : (proc_7_data_FIFO_blk[18] | proc_7_data_PIPO_blk[18] | proc_7_start_FIFO_blk[18] | proc_7_TLF_FIFO_blk[18] | proc_7_input_sync_blk[18] | proc_7_output_sync_blk[18]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_7_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_7_reg <= proc_dep_vld_vec_7;
        end
    end
    assign in_chan_dep_vld_vec_7[0] = dep_chan_vld_0_7;
    assign in_chan_dep_data_vec_7[34 : 0] = dep_chan_data_0_7;
    assign token_in_vec_7[0] = token_0_7;
    assign in_chan_dep_vld_vec_7[1] = dep_chan_vld_1_7;
    assign in_chan_dep_data_vec_7[69 : 35] = dep_chan_data_1_7;
    assign token_in_vec_7[1] = token_1_7;
    assign in_chan_dep_vld_vec_7[2] = dep_chan_vld_2_7;
    assign in_chan_dep_data_vec_7[104 : 70] = dep_chan_data_2_7;
    assign token_in_vec_7[2] = token_2_7;
    assign in_chan_dep_vld_vec_7[3] = dep_chan_vld_3_7;
    assign in_chan_dep_data_vec_7[139 : 105] = dep_chan_data_3_7;
    assign token_in_vec_7[3] = token_3_7;
    assign in_chan_dep_vld_vec_7[4] = dep_chan_vld_4_7;
    assign in_chan_dep_data_vec_7[174 : 140] = dep_chan_data_4_7;
    assign token_in_vec_7[4] = token_4_7;
    assign in_chan_dep_vld_vec_7[5] = dep_chan_vld_5_7;
    assign in_chan_dep_data_vec_7[209 : 175] = dep_chan_data_5_7;
    assign token_in_vec_7[5] = token_5_7;
    assign in_chan_dep_vld_vec_7[6] = dep_chan_vld_6_7;
    assign in_chan_dep_data_vec_7[244 : 210] = dep_chan_data_6_7;
    assign token_in_vec_7[6] = token_6_7;
    assign in_chan_dep_vld_vec_7[7] = dep_chan_vld_8_7;
    assign in_chan_dep_data_vec_7[279 : 245] = dep_chan_data_8_7;
    assign token_in_vec_7[7] = token_8_7;
    assign in_chan_dep_vld_vec_7[8] = dep_chan_vld_9_7;
    assign in_chan_dep_data_vec_7[314 : 280] = dep_chan_data_9_7;
    assign token_in_vec_7[8] = token_9_7;
    assign in_chan_dep_vld_vec_7[9] = dep_chan_vld_10_7;
    assign in_chan_dep_data_vec_7[349 : 315] = dep_chan_data_10_7;
    assign token_in_vec_7[9] = token_10_7;
    assign in_chan_dep_vld_vec_7[10] = dep_chan_vld_11_7;
    assign in_chan_dep_data_vec_7[384 : 350] = dep_chan_data_11_7;
    assign token_in_vec_7[10] = token_11_7;
    assign in_chan_dep_vld_vec_7[11] = dep_chan_vld_12_7;
    assign in_chan_dep_data_vec_7[419 : 385] = dep_chan_data_12_7;
    assign token_in_vec_7[11] = token_12_7;
    assign in_chan_dep_vld_vec_7[12] = dep_chan_vld_13_7;
    assign in_chan_dep_data_vec_7[454 : 420] = dep_chan_data_13_7;
    assign token_in_vec_7[12] = token_13_7;
    assign in_chan_dep_vld_vec_7[13] = dep_chan_vld_14_7;
    assign in_chan_dep_data_vec_7[489 : 455] = dep_chan_data_14_7;
    assign token_in_vec_7[13] = token_14_7;
    assign in_chan_dep_vld_vec_7[14] = dep_chan_vld_15_7;
    assign in_chan_dep_data_vec_7[524 : 490] = dep_chan_data_15_7;
    assign token_in_vec_7[14] = token_15_7;
    assign in_chan_dep_vld_vec_7[15] = dep_chan_vld_16_7;
    assign in_chan_dep_data_vec_7[559 : 525] = dep_chan_data_16_7;
    assign token_in_vec_7[15] = token_16_7;
    assign in_chan_dep_vld_vec_7[16] = dep_chan_vld_17_7;
    assign in_chan_dep_data_vec_7[594 : 560] = dep_chan_data_17_7;
    assign token_in_vec_7[16] = token_17_7;
    assign in_chan_dep_vld_vec_7[17] = dep_chan_vld_18_7;
    assign in_chan_dep_data_vec_7[629 : 595] = dep_chan_data_18_7;
    assign token_in_vec_7[17] = token_18_7;
    assign in_chan_dep_vld_vec_7[18] = dep_chan_vld_23_7;
    assign in_chan_dep_data_vec_7[664 : 630] = dep_chan_data_23_7;
    assign token_in_vec_7[18] = token_23_7;
    assign dep_chan_vld_7_0 = out_chan_dep_vld_vec_7[0];
    assign dep_chan_data_7_0 = out_chan_dep_data_7;
    assign token_7_0 = token_out_vec_7[0];
    assign dep_chan_vld_7_1 = out_chan_dep_vld_vec_7[1];
    assign dep_chan_data_7_1 = out_chan_dep_data_7;
    assign token_7_1 = token_out_vec_7[1];
    assign dep_chan_vld_7_23 = out_chan_dep_vld_vec_7[2];
    assign dep_chan_data_7_23 = out_chan_dep_data_7;
    assign token_7_23 = token_out_vec_7[2];
    assign dep_chan_vld_7_2 = out_chan_dep_vld_vec_7[3];
    assign dep_chan_data_7_2 = out_chan_dep_data_7;
    assign token_7_2 = token_out_vec_7[3];
    assign dep_chan_vld_7_3 = out_chan_dep_vld_vec_7[4];
    assign dep_chan_data_7_3 = out_chan_dep_data_7;
    assign token_7_3 = token_out_vec_7[4];
    assign dep_chan_vld_7_4 = out_chan_dep_vld_vec_7[5];
    assign dep_chan_data_7_4 = out_chan_dep_data_7;
    assign token_7_4 = token_out_vec_7[5];
    assign dep_chan_vld_7_5 = out_chan_dep_vld_vec_7[6];
    assign dep_chan_data_7_5 = out_chan_dep_data_7;
    assign token_7_5 = token_out_vec_7[6];
    assign dep_chan_vld_7_6 = out_chan_dep_vld_vec_7[7];
    assign dep_chan_data_7_6 = out_chan_dep_data_7;
    assign token_7_6 = token_out_vec_7[7];
    assign dep_chan_vld_7_8 = out_chan_dep_vld_vec_7[8];
    assign dep_chan_data_7_8 = out_chan_dep_data_7;
    assign token_7_8 = token_out_vec_7[8];
    assign dep_chan_vld_7_9 = out_chan_dep_vld_vec_7[9];
    assign dep_chan_data_7_9 = out_chan_dep_data_7;
    assign token_7_9 = token_out_vec_7[9];
    assign dep_chan_vld_7_10 = out_chan_dep_vld_vec_7[10];
    assign dep_chan_data_7_10 = out_chan_dep_data_7;
    assign token_7_10 = token_out_vec_7[10];
    assign dep_chan_vld_7_11 = out_chan_dep_vld_vec_7[11];
    assign dep_chan_data_7_11 = out_chan_dep_data_7;
    assign token_7_11 = token_out_vec_7[11];
    assign dep_chan_vld_7_12 = out_chan_dep_vld_vec_7[12];
    assign dep_chan_data_7_12 = out_chan_dep_data_7;
    assign token_7_12 = token_out_vec_7[12];
    assign dep_chan_vld_7_13 = out_chan_dep_vld_vec_7[13];
    assign dep_chan_data_7_13 = out_chan_dep_data_7;
    assign token_7_13 = token_out_vec_7[13];
    assign dep_chan_vld_7_14 = out_chan_dep_vld_vec_7[14];
    assign dep_chan_data_7_14 = out_chan_dep_data_7;
    assign token_7_14 = token_out_vec_7[14];
    assign dep_chan_vld_7_15 = out_chan_dep_vld_vec_7[15];
    assign dep_chan_data_7_15 = out_chan_dep_data_7;
    assign token_7_15 = token_out_vec_7[15];
    assign dep_chan_vld_7_16 = out_chan_dep_vld_vec_7[16];
    assign dep_chan_data_7_16 = out_chan_dep_data_7;
    assign token_7_16 = token_out_vec_7[16];
    assign dep_chan_vld_7_17 = out_chan_dep_vld_vec_7[17];
    assign dep_chan_data_7_17 = out_chan_dep_data_7;
    assign token_7_17 = token_out_vec_7[17];
    assign dep_chan_vld_7_18 = out_chan_dep_vld_vec_7[18];
    assign dep_chan_data_7_18 = out_chan_dep_data_7;
    assign token_7_18 = token_out_vec_7[18];

    // Process: load_value37_U0
    kernel_pr_hls_deadlock_detect_unit #(35, 8, 19, 19) kernel_pr_hls_deadlock_detect_unit_8 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_8),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_8),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_8),
        .token_in_vec(token_in_vec_8),
        .dl_detect_in(dl_detect_out),
        .origin(origin[8]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_8),
        .out_chan_dep_data(out_chan_dep_data_8),
        .token_out_vec(token_out_vec_8),
        .dl_detect_out(dl_in_vec[8]));

    assign proc_8_data_FIFO_blk[0] = 1'b0 | (~load_value37_U0.value_r_blk_n);
    assign proc_8_data_PIPO_blk[0] = 1'b0;
    assign proc_8_start_FIFO_blk[0] = 1'b0;
    assign proc_8_TLF_FIFO_blk[0] = 1'b0;
    assign proc_8_input_sync_blk[0] = 1'b0 | (ap_sync_load_value37_U0_ap_ready & load_value37_U0.ap_idle & ~ap_sync_kernel_pr_entry98_U0_ap_ready);
    assign proc_8_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_8[0] = dl_detect_out ? proc_dep_vld_vec_8_reg[0] : (proc_8_data_FIFO_blk[0] | proc_8_data_PIPO_blk[0] | proc_8_start_FIFO_blk[0] | proc_8_TLF_FIFO_blk[0] | proc_8_input_sync_blk[0] | proc_8_output_sync_blk[0]);
    assign proc_8_data_FIFO_blk[1] = 1'b0 | (~load_value37_U0.bipedge_size_blk_n) | (~load_value37_U0.bipedge_stream_V_V5_blk_n);
    assign proc_8_data_PIPO_blk[1] = 1'b0;
    assign proc_8_start_FIFO_blk[1] = 1'b0;
    assign proc_8_TLF_FIFO_blk[1] = 1'b0;
    assign proc_8_input_sync_blk[1] = 1'b0 | (ap_sync_load_value37_U0_ap_ready & load_value37_U0.ap_idle & ~ap_sync_load_bipedge30_U0_ap_ready);
    assign proc_8_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_8[1] = dl_detect_out ? proc_dep_vld_vec_8_reg[1] : (proc_8_data_FIFO_blk[1] | proc_8_data_PIPO_blk[1] | proc_8_start_FIFO_blk[1] | proc_8_TLF_FIFO_blk[1] | proc_8_input_sync_blk[1] | proc_8_output_sync_blk[1]);
    assign proc_8_data_FIFO_blk[2] = 1'b0 | (~load_value37_U0.value_stream_V_V20_blk_n);
    assign proc_8_data_PIPO_blk[2] = 1'b0;
    assign proc_8_start_FIFO_blk[2] = 1'b0;
    assign proc_8_TLF_FIFO_blk[2] = 1'b0;
    assign proc_8_input_sync_blk[2] = 1'b0;
    assign proc_8_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_8[2] = dl_detect_out ? proc_dep_vld_vec_8_reg[2] : (proc_8_data_FIFO_blk[2] | proc_8_data_PIPO_blk[2] | proc_8_start_FIFO_blk[2] | proc_8_TLF_FIFO_blk[2] | proc_8_input_sync_blk[2] | proc_8_output_sync_blk[2]);
    assign proc_8_data_FIFO_blk[3] = 1'b0;
    assign proc_8_data_PIPO_blk[3] = 1'b0;
    assign proc_8_start_FIFO_blk[3] = 1'b0;
    assign proc_8_TLF_FIFO_blk[3] = 1'b0;
    assign proc_8_input_sync_blk[3] = 1'b0 | (ap_sync_load_value37_U0_ap_ready & load_value37_U0.ap_idle & ~ap_sync_load_bipedge31_U0_ap_ready);
    assign proc_8_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_8[3] = dl_detect_out ? proc_dep_vld_vec_8_reg[3] : (proc_8_data_FIFO_blk[3] | proc_8_data_PIPO_blk[3] | proc_8_start_FIFO_blk[3] | proc_8_TLF_FIFO_blk[3] | proc_8_input_sync_blk[3] | proc_8_output_sync_blk[3]);
    assign proc_8_data_FIFO_blk[4] = 1'b0;
    assign proc_8_data_PIPO_blk[4] = 1'b0;
    assign proc_8_start_FIFO_blk[4] = 1'b0;
    assign proc_8_TLF_FIFO_blk[4] = 1'b0;
    assign proc_8_input_sync_blk[4] = 1'b0 | (ap_sync_load_value37_U0_ap_ready & load_value37_U0.ap_idle & ~ap_sync_load_value32_U0_ap_ready);
    assign proc_8_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_8[4] = dl_detect_out ? proc_dep_vld_vec_8_reg[4] : (proc_8_data_FIFO_blk[4] | proc_8_data_PIPO_blk[4] | proc_8_start_FIFO_blk[4] | proc_8_TLF_FIFO_blk[4] | proc_8_input_sync_blk[4] | proc_8_output_sync_blk[4]);
    assign proc_8_data_FIFO_blk[5] = 1'b0;
    assign proc_8_data_PIPO_blk[5] = 1'b0;
    assign proc_8_start_FIFO_blk[5] = 1'b0;
    assign proc_8_TLF_FIFO_blk[5] = 1'b0;
    assign proc_8_input_sync_blk[5] = 1'b0 | (ap_sync_load_value37_U0_ap_ready & load_value37_U0.ap_idle & ~ap_sync_load_value33_U0_ap_ready);
    assign proc_8_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_8[5] = dl_detect_out ? proc_dep_vld_vec_8_reg[5] : (proc_8_data_FIFO_blk[5] | proc_8_data_PIPO_blk[5] | proc_8_start_FIFO_blk[5] | proc_8_TLF_FIFO_blk[5] | proc_8_input_sync_blk[5] | proc_8_output_sync_blk[5]);
    assign proc_8_data_FIFO_blk[6] = 1'b0;
    assign proc_8_data_PIPO_blk[6] = 1'b0;
    assign proc_8_start_FIFO_blk[6] = 1'b0;
    assign proc_8_TLF_FIFO_blk[6] = 1'b0;
    assign proc_8_input_sync_blk[6] = 1'b0 | (ap_sync_load_value37_U0_ap_ready & load_value37_U0.ap_idle & ~ap_sync_load_value34_U0_ap_ready);
    assign proc_8_output_sync_blk[6] = 1'b0;
    assign proc_dep_vld_vec_8[6] = dl_detect_out ? proc_dep_vld_vec_8_reg[6] : (proc_8_data_FIFO_blk[6] | proc_8_data_PIPO_blk[6] | proc_8_start_FIFO_blk[6] | proc_8_TLF_FIFO_blk[6] | proc_8_input_sync_blk[6] | proc_8_output_sync_blk[6]);
    assign proc_8_data_FIFO_blk[7] = 1'b0;
    assign proc_8_data_PIPO_blk[7] = 1'b0;
    assign proc_8_start_FIFO_blk[7] = 1'b0;
    assign proc_8_TLF_FIFO_blk[7] = 1'b0;
    assign proc_8_input_sync_blk[7] = 1'b0 | (ap_sync_load_value37_U0_ap_ready & load_value37_U0.ap_idle & ~ap_sync_load_value35_U0_ap_ready);
    assign proc_8_output_sync_blk[7] = 1'b0;
    assign proc_dep_vld_vec_8[7] = dl_detect_out ? proc_dep_vld_vec_8_reg[7] : (proc_8_data_FIFO_blk[7] | proc_8_data_PIPO_blk[7] | proc_8_start_FIFO_blk[7] | proc_8_TLF_FIFO_blk[7] | proc_8_input_sync_blk[7] | proc_8_output_sync_blk[7]);
    assign proc_8_data_FIFO_blk[8] = 1'b0;
    assign proc_8_data_PIPO_blk[8] = 1'b0;
    assign proc_8_start_FIFO_blk[8] = 1'b0;
    assign proc_8_TLF_FIFO_blk[8] = 1'b0;
    assign proc_8_input_sync_blk[8] = 1'b0 | (ap_sync_load_value37_U0_ap_ready & load_value37_U0.ap_idle & ~ap_sync_load_value36_U0_ap_ready);
    assign proc_8_output_sync_blk[8] = 1'b0;
    assign proc_dep_vld_vec_8[8] = dl_detect_out ? proc_dep_vld_vec_8_reg[8] : (proc_8_data_FIFO_blk[8] | proc_8_data_PIPO_blk[8] | proc_8_start_FIFO_blk[8] | proc_8_TLF_FIFO_blk[8] | proc_8_input_sync_blk[8] | proc_8_output_sync_blk[8]);
    assign proc_8_data_FIFO_blk[9] = 1'b0;
    assign proc_8_data_PIPO_blk[9] = 1'b0;
    assign proc_8_start_FIFO_blk[9] = 1'b0;
    assign proc_8_TLF_FIFO_blk[9] = 1'b0;
    assign proc_8_input_sync_blk[9] = 1'b0 | (ap_sync_load_value37_U0_ap_ready & load_value37_U0.ap_idle & ~ap_sync_load_value38_U0_ap_ready);
    assign proc_8_output_sync_blk[9] = 1'b0;
    assign proc_dep_vld_vec_8[9] = dl_detect_out ? proc_dep_vld_vec_8_reg[9] : (proc_8_data_FIFO_blk[9] | proc_8_data_PIPO_blk[9] | proc_8_start_FIFO_blk[9] | proc_8_TLF_FIFO_blk[9] | proc_8_input_sync_blk[9] | proc_8_output_sync_blk[9]);
    assign proc_8_data_FIFO_blk[10] = 1'b0;
    assign proc_8_data_PIPO_blk[10] = 1'b0;
    assign proc_8_start_FIFO_blk[10] = 1'b0;
    assign proc_8_TLF_FIFO_blk[10] = 1'b0;
    assign proc_8_input_sync_blk[10] = 1'b0 | (ap_sync_load_value37_U0_ap_ready & load_value37_U0.ap_idle & ~ap_sync_load_value39_U0_ap_ready);
    assign proc_8_output_sync_blk[10] = 1'b0;
    assign proc_dep_vld_vec_8[10] = dl_detect_out ? proc_dep_vld_vec_8_reg[10] : (proc_8_data_FIFO_blk[10] | proc_8_data_PIPO_blk[10] | proc_8_start_FIFO_blk[10] | proc_8_TLF_FIFO_blk[10] | proc_8_input_sync_blk[10] | proc_8_output_sync_blk[10]);
    assign proc_8_data_FIFO_blk[11] = 1'b0;
    assign proc_8_data_PIPO_blk[11] = 1'b0;
    assign proc_8_start_FIFO_blk[11] = 1'b0;
    assign proc_8_TLF_FIFO_blk[11] = 1'b0;
    assign proc_8_input_sync_blk[11] = 1'b0 | (ap_sync_load_value37_U0_ap_ready & load_value37_U0.ap_idle & ~ap_sync_load_value40_U0_ap_ready);
    assign proc_8_output_sync_blk[11] = 1'b0;
    assign proc_dep_vld_vec_8[11] = dl_detect_out ? proc_dep_vld_vec_8_reg[11] : (proc_8_data_FIFO_blk[11] | proc_8_data_PIPO_blk[11] | proc_8_start_FIFO_blk[11] | proc_8_TLF_FIFO_blk[11] | proc_8_input_sync_blk[11] | proc_8_output_sync_blk[11]);
    assign proc_8_data_FIFO_blk[12] = 1'b0;
    assign proc_8_data_PIPO_blk[12] = 1'b0;
    assign proc_8_start_FIFO_blk[12] = 1'b0;
    assign proc_8_TLF_FIFO_blk[12] = 1'b0;
    assign proc_8_input_sync_blk[12] = 1'b0 | (ap_sync_load_value37_U0_ap_ready & load_value37_U0.ap_idle & ~ap_sync_load_value41_U0_ap_ready);
    assign proc_8_output_sync_blk[12] = 1'b0;
    assign proc_dep_vld_vec_8[12] = dl_detect_out ? proc_dep_vld_vec_8_reg[12] : (proc_8_data_FIFO_blk[12] | proc_8_data_PIPO_blk[12] | proc_8_start_FIFO_blk[12] | proc_8_TLF_FIFO_blk[12] | proc_8_input_sync_blk[12] | proc_8_output_sync_blk[12]);
    assign proc_8_data_FIFO_blk[13] = 1'b0;
    assign proc_8_data_PIPO_blk[13] = 1'b0;
    assign proc_8_start_FIFO_blk[13] = 1'b0;
    assign proc_8_TLF_FIFO_blk[13] = 1'b0;
    assign proc_8_input_sync_blk[13] = 1'b0 | (ap_sync_load_value37_U0_ap_ready & load_value37_U0.ap_idle & ~ap_sync_load_value42_U0_ap_ready);
    assign proc_8_output_sync_blk[13] = 1'b0;
    assign proc_dep_vld_vec_8[13] = dl_detect_out ? proc_dep_vld_vec_8_reg[13] : (proc_8_data_FIFO_blk[13] | proc_8_data_PIPO_blk[13] | proc_8_start_FIFO_blk[13] | proc_8_TLF_FIFO_blk[13] | proc_8_input_sync_blk[13] | proc_8_output_sync_blk[13]);
    assign proc_8_data_FIFO_blk[14] = 1'b0;
    assign proc_8_data_PIPO_blk[14] = 1'b0;
    assign proc_8_start_FIFO_blk[14] = 1'b0;
    assign proc_8_TLF_FIFO_blk[14] = 1'b0;
    assign proc_8_input_sync_blk[14] = 1'b0 | (ap_sync_load_value37_U0_ap_ready & load_value37_U0.ap_idle & ~ap_sync_load_value43_U0_ap_ready);
    assign proc_8_output_sync_blk[14] = 1'b0;
    assign proc_dep_vld_vec_8[14] = dl_detect_out ? proc_dep_vld_vec_8_reg[14] : (proc_8_data_FIFO_blk[14] | proc_8_data_PIPO_blk[14] | proc_8_start_FIFO_blk[14] | proc_8_TLF_FIFO_blk[14] | proc_8_input_sync_blk[14] | proc_8_output_sync_blk[14]);
    assign proc_8_data_FIFO_blk[15] = 1'b0;
    assign proc_8_data_PIPO_blk[15] = 1'b0;
    assign proc_8_start_FIFO_blk[15] = 1'b0;
    assign proc_8_TLF_FIFO_blk[15] = 1'b0;
    assign proc_8_input_sync_blk[15] = 1'b0 | (ap_sync_load_value37_U0_ap_ready & load_value37_U0.ap_idle & ~ap_sync_load_value44_U0_ap_ready);
    assign proc_8_output_sync_blk[15] = 1'b0;
    assign proc_dep_vld_vec_8[15] = dl_detect_out ? proc_dep_vld_vec_8_reg[15] : (proc_8_data_FIFO_blk[15] | proc_8_data_PIPO_blk[15] | proc_8_start_FIFO_blk[15] | proc_8_TLF_FIFO_blk[15] | proc_8_input_sync_blk[15] | proc_8_output_sync_blk[15]);
    assign proc_8_data_FIFO_blk[16] = 1'b0;
    assign proc_8_data_PIPO_blk[16] = 1'b0;
    assign proc_8_start_FIFO_blk[16] = 1'b0;
    assign proc_8_TLF_FIFO_blk[16] = 1'b0;
    assign proc_8_input_sync_blk[16] = 1'b0 | (ap_sync_load_value37_U0_ap_ready & load_value37_U0.ap_idle & ~ap_sync_load_value45_U0_ap_ready);
    assign proc_8_output_sync_blk[16] = 1'b0;
    assign proc_dep_vld_vec_8[16] = dl_detect_out ? proc_dep_vld_vec_8_reg[16] : (proc_8_data_FIFO_blk[16] | proc_8_data_PIPO_blk[16] | proc_8_start_FIFO_blk[16] | proc_8_TLF_FIFO_blk[16] | proc_8_input_sync_blk[16] | proc_8_output_sync_blk[16]);
    assign proc_8_data_FIFO_blk[17] = 1'b0;
    assign proc_8_data_PIPO_blk[17] = 1'b0;
    assign proc_8_start_FIFO_blk[17] = 1'b0;
    assign proc_8_TLF_FIFO_blk[17] = 1'b0;
    assign proc_8_input_sync_blk[17] = 1'b0 | (ap_sync_load_value37_U0_ap_ready & load_value37_U0.ap_idle & ~ap_sync_load_value46_U0_ap_ready);
    assign proc_8_output_sync_blk[17] = 1'b0;
    assign proc_dep_vld_vec_8[17] = dl_detect_out ? proc_dep_vld_vec_8_reg[17] : (proc_8_data_FIFO_blk[17] | proc_8_data_PIPO_blk[17] | proc_8_start_FIFO_blk[17] | proc_8_TLF_FIFO_blk[17] | proc_8_input_sync_blk[17] | proc_8_output_sync_blk[17]);
    assign proc_8_data_FIFO_blk[18] = 1'b0;
    assign proc_8_data_PIPO_blk[18] = 1'b0;
    assign proc_8_start_FIFO_blk[18] = 1'b0;
    assign proc_8_TLF_FIFO_blk[18] = 1'b0;
    assign proc_8_input_sync_blk[18] = 1'b0 | (ap_sync_load_value37_U0_ap_ready & load_value37_U0.ap_idle & ~ap_sync_load_value47_U0_ap_ready);
    assign proc_8_output_sync_blk[18] = 1'b0;
    assign proc_dep_vld_vec_8[18] = dl_detect_out ? proc_dep_vld_vec_8_reg[18] : (proc_8_data_FIFO_blk[18] | proc_8_data_PIPO_blk[18] | proc_8_start_FIFO_blk[18] | proc_8_TLF_FIFO_blk[18] | proc_8_input_sync_blk[18] | proc_8_output_sync_blk[18]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_8_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_8_reg <= proc_dep_vld_vec_8;
        end
    end
    assign in_chan_dep_vld_vec_8[0] = dep_chan_vld_0_8;
    assign in_chan_dep_data_vec_8[34 : 0] = dep_chan_data_0_8;
    assign token_in_vec_8[0] = token_0_8;
    assign in_chan_dep_vld_vec_8[1] = dep_chan_vld_1_8;
    assign in_chan_dep_data_vec_8[69 : 35] = dep_chan_data_1_8;
    assign token_in_vec_8[1] = token_1_8;
    assign in_chan_dep_vld_vec_8[2] = dep_chan_vld_2_8;
    assign in_chan_dep_data_vec_8[104 : 70] = dep_chan_data_2_8;
    assign token_in_vec_8[2] = token_2_8;
    assign in_chan_dep_vld_vec_8[3] = dep_chan_vld_3_8;
    assign in_chan_dep_data_vec_8[139 : 105] = dep_chan_data_3_8;
    assign token_in_vec_8[3] = token_3_8;
    assign in_chan_dep_vld_vec_8[4] = dep_chan_vld_4_8;
    assign in_chan_dep_data_vec_8[174 : 140] = dep_chan_data_4_8;
    assign token_in_vec_8[4] = token_4_8;
    assign in_chan_dep_vld_vec_8[5] = dep_chan_vld_5_8;
    assign in_chan_dep_data_vec_8[209 : 175] = dep_chan_data_5_8;
    assign token_in_vec_8[5] = token_5_8;
    assign in_chan_dep_vld_vec_8[6] = dep_chan_vld_6_8;
    assign in_chan_dep_data_vec_8[244 : 210] = dep_chan_data_6_8;
    assign token_in_vec_8[6] = token_6_8;
    assign in_chan_dep_vld_vec_8[7] = dep_chan_vld_7_8;
    assign in_chan_dep_data_vec_8[279 : 245] = dep_chan_data_7_8;
    assign token_in_vec_8[7] = token_7_8;
    assign in_chan_dep_vld_vec_8[8] = dep_chan_vld_9_8;
    assign in_chan_dep_data_vec_8[314 : 280] = dep_chan_data_9_8;
    assign token_in_vec_8[8] = token_9_8;
    assign in_chan_dep_vld_vec_8[9] = dep_chan_vld_10_8;
    assign in_chan_dep_data_vec_8[349 : 315] = dep_chan_data_10_8;
    assign token_in_vec_8[9] = token_10_8;
    assign in_chan_dep_vld_vec_8[10] = dep_chan_vld_11_8;
    assign in_chan_dep_data_vec_8[384 : 350] = dep_chan_data_11_8;
    assign token_in_vec_8[10] = token_11_8;
    assign in_chan_dep_vld_vec_8[11] = dep_chan_vld_12_8;
    assign in_chan_dep_data_vec_8[419 : 385] = dep_chan_data_12_8;
    assign token_in_vec_8[11] = token_12_8;
    assign in_chan_dep_vld_vec_8[12] = dep_chan_vld_13_8;
    assign in_chan_dep_data_vec_8[454 : 420] = dep_chan_data_13_8;
    assign token_in_vec_8[12] = token_13_8;
    assign in_chan_dep_vld_vec_8[13] = dep_chan_vld_14_8;
    assign in_chan_dep_data_vec_8[489 : 455] = dep_chan_data_14_8;
    assign token_in_vec_8[13] = token_14_8;
    assign in_chan_dep_vld_vec_8[14] = dep_chan_vld_15_8;
    assign in_chan_dep_data_vec_8[524 : 490] = dep_chan_data_15_8;
    assign token_in_vec_8[14] = token_15_8;
    assign in_chan_dep_vld_vec_8[15] = dep_chan_vld_16_8;
    assign in_chan_dep_data_vec_8[559 : 525] = dep_chan_data_16_8;
    assign token_in_vec_8[15] = token_16_8;
    assign in_chan_dep_vld_vec_8[16] = dep_chan_vld_17_8;
    assign in_chan_dep_data_vec_8[594 : 560] = dep_chan_data_17_8;
    assign token_in_vec_8[16] = token_17_8;
    assign in_chan_dep_vld_vec_8[17] = dep_chan_vld_18_8;
    assign in_chan_dep_data_vec_8[629 : 595] = dep_chan_data_18_8;
    assign token_in_vec_8[17] = token_18_8;
    assign in_chan_dep_vld_vec_8[18] = dep_chan_vld_24_8;
    assign in_chan_dep_data_vec_8[664 : 630] = dep_chan_data_24_8;
    assign token_in_vec_8[18] = token_24_8;
    assign dep_chan_vld_8_0 = out_chan_dep_vld_vec_8[0];
    assign dep_chan_data_8_0 = out_chan_dep_data_8;
    assign token_8_0 = token_out_vec_8[0];
    assign dep_chan_vld_8_1 = out_chan_dep_vld_vec_8[1];
    assign dep_chan_data_8_1 = out_chan_dep_data_8;
    assign token_8_1 = token_out_vec_8[1];
    assign dep_chan_vld_8_24 = out_chan_dep_vld_vec_8[2];
    assign dep_chan_data_8_24 = out_chan_dep_data_8;
    assign token_8_24 = token_out_vec_8[2];
    assign dep_chan_vld_8_2 = out_chan_dep_vld_vec_8[3];
    assign dep_chan_data_8_2 = out_chan_dep_data_8;
    assign token_8_2 = token_out_vec_8[3];
    assign dep_chan_vld_8_3 = out_chan_dep_vld_vec_8[4];
    assign dep_chan_data_8_3 = out_chan_dep_data_8;
    assign token_8_3 = token_out_vec_8[4];
    assign dep_chan_vld_8_4 = out_chan_dep_vld_vec_8[5];
    assign dep_chan_data_8_4 = out_chan_dep_data_8;
    assign token_8_4 = token_out_vec_8[5];
    assign dep_chan_vld_8_5 = out_chan_dep_vld_vec_8[6];
    assign dep_chan_data_8_5 = out_chan_dep_data_8;
    assign token_8_5 = token_out_vec_8[6];
    assign dep_chan_vld_8_6 = out_chan_dep_vld_vec_8[7];
    assign dep_chan_data_8_6 = out_chan_dep_data_8;
    assign token_8_6 = token_out_vec_8[7];
    assign dep_chan_vld_8_7 = out_chan_dep_vld_vec_8[8];
    assign dep_chan_data_8_7 = out_chan_dep_data_8;
    assign token_8_7 = token_out_vec_8[8];
    assign dep_chan_vld_8_9 = out_chan_dep_vld_vec_8[9];
    assign dep_chan_data_8_9 = out_chan_dep_data_8;
    assign token_8_9 = token_out_vec_8[9];
    assign dep_chan_vld_8_10 = out_chan_dep_vld_vec_8[10];
    assign dep_chan_data_8_10 = out_chan_dep_data_8;
    assign token_8_10 = token_out_vec_8[10];
    assign dep_chan_vld_8_11 = out_chan_dep_vld_vec_8[11];
    assign dep_chan_data_8_11 = out_chan_dep_data_8;
    assign token_8_11 = token_out_vec_8[11];
    assign dep_chan_vld_8_12 = out_chan_dep_vld_vec_8[12];
    assign dep_chan_data_8_12 = out_chan_dep_data_8;
    assign token_8_12 = token_out_vec_8[12];
    assign dep_chan_vld_8_13 = out_chan_dep_vld_vec_8[13];
    assign dep_chan_data_8_13 = out_chan_dep_data_8;
    assign token_8_13 = token_out_vec_8[13];
    assign dep_chan_vld_8_14 = out_chan_dep_vld_vec_8[14];
    assign dep_chan_data_8_14 = out_chan_dep_data_8;
    assign token_8_14 = token_out_vec_8[14];
    assign dep_chan_vld_8_15 = out_chan_dep_vld_vec_8[15];
    assign dep_chan_data_8_15 = out_chan_dep_data_8;
    assign token_8_15 = token_out_vec_8[15];
    assign dep_chan_vld_8_16 = out_chan_dep_vld_vec_8[16];
    assign dep_chan_data_8_16 = out_chan_dep_data_8;
    assign token_8_16 = token_out_vec_8[16];
    assign dep_chan_vld_8_17 = out_chan_dep_vld_vec_8[17];
    assign dep_chan_data_8_17 = out_chan_dep_data_8;
    assign token_8_17 = token_out_vec_8[17];
    assign dep_chan_vld_8_18 = out_chan_dep_vld_vec_8[18];
    assign dep_chan_data_8_18 = out_chan_dep_data_8;
    assign token_8_18 = token_out_vec_8[18];

    // Process: load_value38_U0
    kernel_pr_hls_deadlock_detect_unit #(35, 9, 19, 19) kernel_pr_hls_deadlock_detect_unit_9 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_9),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_9),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_9),
        .token_in_vec(token_in_vec_9),
        .dl_detect_in(dl_detect_out),
        .origin(origin[9]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_9),
        .out_chan_dep_data(out_chan_dep_data_9),
        .token_out_vec(token_out_vec_9),
        .dl_detect_out(dl_in_vec[9]));

    assign proc_9_data_FIFO_blk[0] = 1'b0 | (~load_value38_U0.value_r_blk_n);
    assign proc_9_data_PIPO_blk[0] = 1'b0;
    assign proc_9_start_FIFO_blk[0] = 1'b0;
    assign proc_9_TLF_FIFO_blk[0] = 1'b0;
    assign proc_9_input_sync_blk[0] = 1'b0 | (ap_sync_load_value38_U0_ap_ready & load_value38_U0.ap_idle & ~ap_sync_kernel_pr_entry98_U0_ap_ready);
    assign proc_9_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_9[0] = dl_detect_out ? proc_dep_vld_vec_9_reg[0] : (proc_9_data_FIFO_blk[0] | proc_9_data_PIPO_blk[0] | proc_9_start_FIFO_blk[0] | proc_9_TLF_FIFO_blk[0] | proc_9_input_sync_blk[0] | proc_9_output_sync_blk[0]);
    assign proc_9_data_FIFO_blk[1] = 1'b0 | (~load_value38_U0.bipedge_size_blk_n) | (~load_value38_U0.bipedge_stream_V_V6_blk_n);
    assign proc_9_data_PIPO_blk[1] = 1'b0;
    assign proc_9_start_FIFO_blk[1] = 1'b0;
    assign proc_9_TLF_FIFO_blk[1] = 1'b0;
    assign proc_9_input_sync_blk[1] = 1'b0 | (ap_sync_load_value38_U0_ap_ready & load_value38_U0.ap_idle & ~ap_sync_load_bipedge30_U0_ap_ready);
    assign proc_9_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_9[1] = dl_detect_out ? proc_dep_vld_vec_9_reg[1] : (proc_9_data_FIFO_blk[1] | proc_9_data_PIPO_blk[1] | proc_9_start_FIFO_blk[1] | proc_9_TLF_FIFO_blk[1] | proc_9_input_sync_blk[1] | proc_9_output_sync_blk[1]);
    assign proc_9_data_FIFO_blk[2] = 1'b0 | (~load_value38_U0.value_stream_V_V21_blk_n);
    assign proc_9_data_PIPO_blk[2] = 1'b0;
    assign proc_9_start_FIFO_blk[2] = 1'b0;
    assign proc_9_TLF_FIFO_blk[2] = 1'b0;
    assign proc_9_input_sync_blk[2] = 1'b0;
    assign proc_9_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_9[2] = dl_detect_out ? proc_dep_vld_vec_9_reg[2] : (proc_9_data_FIFO_blk[2] | proc_9_data_PIPO_blk[2] | proc_9_start_FIFO_blk[2] | proc_9_TLF_FIFO_blk[2] | proc_9_input_sync_blk[2] | proc_9_output_sync_blk[2]);
    assign proc_9_data_FIFO_blk[3] = 1'b0;
    assign proc_9_data_PIPO_blk[3] = 1'b0;
    assign proc_9_start_FIFO_blk[3] = 1'b0;
    assign proc_9_TLF_FIFO_blk[3] = 1'b0;
    assign proc_9_input_sync_blk[3] = 1'b0 | (ap_sync_load_value38_U0_ap_ready & load_value38_U0.ap_idle & ~ap_sync_load_bipedge31_U0_ap_ready);
    assign proc_9_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_9[3] = dl_detect_out ? proc_dep_vld_vec_9_reg[3] : (proc_9_data_FIFO_blk[3] | proc_9_data_PIPO_blk[3] | proc_9_start_FIFO_blk[3] | proc_9_TLF_FIFO_blk[3] | proc_9_input_sync_blk[3] | proc_9_output_sync_blk[3]);
    assign proc_9_data_FIFO_blk[4] = 1'b0;
    assign proc_9_data_PIPO_blk[4] = 1'b0;
    assign proc_9_start_FIFO_blk[4] = 1'b0;
    assign proc_9_TLF_FIFO_blk[4] = 1'b0;
    assign proc_9_input_sync_blk[4] = 1'b0 | (ap_sync_load_value38_U0_ap_ready & load_value38_U0.ap_idle & ~ap_sync_load_value32_U0_ap_ready);
    assign proc_9_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_9[4] = dl_detect_out ? proc_dep_vld_vec_9_reg[4] : (proc_9_data_FIFO_blk[4] | proc_9_data_PIPO_blk[4] | proc_9_start_FIFO_blk[4] | proc_9_TLF_FIFO_blk[4] | proc_9_input_sync_blk[4] | proc_9_output_sync_blk[4]);
    assign proc_9_data_FIFO_blk[5] = 1'b0;
    assign proc_9_data_PIPO_blk[5] = 1'b0;
    assign proc_9_start_FIFO_blk[5] = 1'b0;
    assign proc_9_TLF_FIFO_blk[5] = 1'b0;
    assign proc_9_input_sync_blk[5] = 1'b0 | (ap_sync_load_value38_U0_ap_ready & load_value38_U0.ap_idle & ~ap_sync_load_value33_U0_ap_ready);
    assign proc_9_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_9[5] = dl_detect_out ? proc_dep_vld_vec_9_reg[5] : (proc_9_data_FIFO_blk[5] | proc_9_data_PIPO_blk[5] | proc_9_start_FIFO_blk[5] | proc_9_TLF_FIFO_blk[5] | proc_9_input_sync_blk[5] | proc_9_output_sync_blk[5]);
    assign proc_9_data_FIFO_blk[6] = 1'b0;
    assign proc_9_data_PIPO_blk[6] = 1'b0;
    assign proc_9_start_FIFO_blk[6] = 1'b0;
    assign proc_9_TLF_FIFO_blk[6] = 1'b0;
    assign proc_9_input_sync_blk[6] = 1'b0 | (ap_sync_load_value38_U0_ap_ready & load_value38_U0.ap_idle & ~ap_sync_load_value34_U0_ap_ready);
    assign proc_9_output_sync_blk[6] = 1'b0;
    assign proc_dep_vld_vec_9[6] = dl_detect_out ? proc_dep_vld_vec_9_reg[6] : (proc_9_data_FIFO_blk[6] | proc_9_data_PIPO_blk[6] | proc_9_start_FIFO_blk[6] | proc_9_TLF_FIFO_blk[6] | proc_9_input_sync_blk[6] | proc_9_output_sync_blk[6]);
    assign proc_9_data_FIFO_blk[7] = 1'b0;
    assign proc_9_data_PIPO_blk[7] = 1'b0;
    assign proc_9_start_FIFO_blk[7] = 1'b0;
    assign proc_9_TLF_FIFO_blk[7] = 1'b0;
    assign proc_9_input_sync_blk[7] = 1'b0 | (ap_sync_load_value38_U0_ap_ready & load_value38_U0.ap_idle & ~ap_sync_load_value35_U0_ap_ready);
    assign proc_9_output_sync_blk[7] = 1'b0;
    assign proc_dep_vld_vec_9[7] = dl_detect_out ? proc_dep_vld_vec_9_reg[7] : (proc_9_data_FIFO_blk[7] | proc_9_data_PIPO_blk[7] | proc_9_start_FIFO_blk[7] | proc_9_TLF_FIFO_blk[7] | proc_9_input_sync_blk[7] | proc_9_output_sync_blk[7]);
    assign proc_9_data_FIFO_blk[8] = 1'b0;
    assign proc_9_data_PIPO_blk[8] = 1'b0;
    assign proc_9_start_FIFO_blk[8] = 1'b0;
    assign proc_9_TLF_FIFO_blk[8] = 1'b0;
    assign proc_9_input_sync_blk[8] = 1'b0 | (ap_sync_load_value38_U0_ap_ready & load_value38_U0.ap_idle & ~ap_sync_load_value36_U0_ap_ready);
    assign proc_9_output_sync_blk[8] = 1'b0;
    assign proc_dep_vld_vec_9[8] = dl_detect_out ? proc_dep_vld_vec_9_reg[8] : (proc_9_data_FIFO_blk[8] | proc_9_data_PIPO_blk[8] | proc_9_start_FIFO_blk[8] | proc_9_TLF_FIFO_blk[8] | proc_9_input_sync_blk[8] | proc_9_output_sync_blk[8]);
    assign proc_9_data_FIFO_blk[9] = 1'b0;
    assign proc_9_data_PIPO_blk[9] = 1'b0;
    assign proc_9_start_FIFO_blk[9] = 1'b0;
    assign proc_9_TLF_FIFO_blk[9] = 1'b0;
    assign proc_9_input_sync_blk[9] = 1'b0 | (ap_sync_load_value38_U0_ap_ready & load_value38_U0.ap_idle & ~ap_sync_load_value37_U0_ap_ready);
    assign proc_9_output_sync_blk[9] = 1'b0;
    assign proc_dep_vld_vec_9[9] = dl_detect_out ? proc_dep_vld_vec_9_reg[9] : (proc_9_data_FIFO_blk[9] | proc_9_data_PIPO_blk[9] | proc_9_start_FIFO_blk[9] | proc_9_TLF_FIFO_blk[9] | proc_9_input_sync_blk[9] | proc_9_output_sync_blk[9]);
    assign proc_9_data_FIFO_blk[10] = 1'b0;
    assign proc_9_data_PIPO_blk[10] = 1'b0;
    assign proc_9_start_FIFO_blk[10] = 1'b0;
    assign proc_9_TLF_FIFO_blk[10] = 1'b0;
    assign proc_9_input_sync_blk[10] = 1'b0 | (ap_sync_load_value38_U0_ap_ready & load_value38_U0.ap_idle & ~ap_sync_load_value39_U0_ap_ready);
    assign proc_9_output_sync_blk[10] = 1'b0;
    assign proc_dep_vld_vec_9[10] = dl_detect_out ? proc_dep_vld_vec_9_reg[10] : (proc_9_data_FIFO_blk[10] | proc_9_data_PIPO_blk[10] | proc_9_start_FIFO_blk[10] | proc_9_TLF_FIFO_blk[10] | proc_9_input_sync_blk[10] | proc_9_output_sync_blk[10]);
    assign proc_9_data_FIFO_blk[11] = 1'b0;
    assign proc_9_data_PIPO_blk[11] = 1'b0;
    assign proc_9_start_FIFO_blk[11] = 1'b0;
    assign proc_9_TLF_FIFO_blk[11] = 1'b0;
    assign proc_9_input_sync_blk[11] = 1'b0 | (ap_sync_load_value38_U0_ap_ready & load_value38_U0.ap_idle & ~ap_sync_load_value40_U0_ap_ready);
    assign proc_9_output_sync_blk[11] = 1'b0;
    assign proc_dep_vld_vec_9[11] = dl_detect_out ? proc_dep_vld_vec_9_reg[11] : (proc_9_data_FIFO_blk[11] | proc_9_data_PIPO_blk[11] | proc_9_start_FIFO_blk[11] | proc_9_TLF_FIFO_blk[11] | proc_9_input_sync_blk[11] | proc_9_output_sync_blk[11]);
    assign proc_9_data_FIFO_blk[12] = 1'b0;
    assign proc_9_data_PIPO_blk[12] = 1'b0;
    assign proc_9_start_FIFO_blk[12] = 1'b0;
    assign proc_9_TLF_FIFO_blk[12] = 1'b0;
    assign proc_9_input_sync_blk[12] = 1'b0 | (ap_sync_load_value38_U0_ap_ready & load_value38_U0.ap_idle & ~ap_sync_load_value41_U0_ap_ready);
    assign proc_9_output_sync_blk[12] = 1'b0;
    assign proc_dep_vld_vec_9[12] = dl_detect_out ? proc_dep_vld_vec_9_reg[12] : (proc_9_data_FIFO_blk[12] | proc_9_data_PIPO_blk[12] | proc_9_start_FIFO_blk[12] | proc_9_TLF_FIFO_blk[12] | proc_9_input_sync_blk[12] | proc_9_output_sync_blk[12]);
    assign proc_9_data_FIFO_blk[13] = 1'b0;
    assign proc_9_data_PIPO_blk[13] = 1'b0;
    assign proc_9_start_FIFO_blk[13] = 1'b0;
    assign proc_9_TLF_FIFO_blk[13] = 1'b0;
    assign proc_9_input_sync_blk[13] = 1'b0 | (ap_sync_load_value38_U0_ap_ready & load_value38_U0.ap_idle & ~ap_sync_load_value42_U0_ap_ready);
    assign proc_9_output_sync_blk[13] = 1'b0;
    assign proc_dep_vld_vec_9[13] = dl_detect_out ? proc_dep_vld_vec_9_reg[13] : (proc_9_data_FIFO_blk[13] | proc_9_data_PIPO_blk[13] | proc_9_start_FIFO_blk[13] | proc_9_TLF_FIFO_blk[13] | proc_9_input_sync_blk[13] | proc_9_output_sync_blk[13]);
    assign proc_9_data_FIFO_blk[14] = 1'b0;
    assign proc_9_data_PIPO_blk[14] = 1'b0;
    assign proc_9_start_FIFO_blk[14] = 1'b0;
    assign proc_9_TLF_FIFO_blk[14] = 1'b0;
    assign proc_9_input_sync_blk[14] = 1'b0 | (ap_sync_load_value38_U0_ap_ready & load_value38_U0.ap_idle & ~ap_sync_load_value43_U0_ap_ready);
    assign proc_9_output_sync_blk[14] = 1'b0;
    assign proc_dep_vld_vec_9[14] = dl_detect_out ? proc_dep_vld_vec_9_reg[14] : (proc_9_data_FIFO_blk[14] | proc_9_data_PIPO_blk[14] | proc_9_start_FIFO_blk[14] | proc_9_TLF_FIFO_blk[14] | proc_9_input_sync_blk[14] | proc_9_output_sync_blk[14]);
    assign proc_9_data_FIFO_blk[15] = 1'b0;
    assign proc_9_data_PIPO_blk[15] = 1'b0;
    assign proc_9_start_FIFO_blk[15] = 1'b0;
    assign proc_9_TLF_FIFO_blk[15] = 1'b0;
    assign proc_9_input_sync_blk[15] = 1'b0 | (ap_sync_load_value38_U0_ap_ready & load_value38_U0.ap_idle & ~ap_sync_load_value44_U0_ap_ready);
    assign proc_9_output_sync_blk[15] = 1'b0;
    assign proc_dep_vld_vec_9[15] = dl_detect_out ? proc_dep_vld_vec_9_reg[15] : (proc_9_data_FIFO_blk[15] | proc_9_data_PIPO_blk[15] | proc_9_start_FIFO_blk[15] | proc_9_TLF_FIFO_blk[15] | proc_9_input_sync_blk[15] | proc_9_output_sync_blk[15]);
    assign proc_9_data_FIFO_blk[16] = 1'b0;
    assign proc_9_data_PIPO_blk[16] = 1'b0;
    assign proc_9_start_FIFO_blk[16] = 1'b0;
    assign proc_9_TLF_FIFO_blk[16] = 1'b0;
    assign proc_9_input_sync_blk[16] = 1'b0 | (ap_sync_load_value38_U0_ap_ready & load_value38_U0.ap_idle & ~ap_sync_load_value45_U0_ap_ready);
    assign proc_9_output_sync_blk[16] = 1'b0;
    assign proc_dep_vld_vec_9[16] = dl_detect_out ? proc_dep_vld_vec_9_reg[16] : (proc_9_data_FIFO_blk[16] | proc_9_data_PIPO_blk[16] | proc_9_start_FIFO_blk[16] | proc_9_TLF_FIFO_blk[16] | proc_9_input_sync_blk[16] | proc_9_output_sync_blk[16]);
    assign proc_9_data_FIFO_blk[17] = 1'b0;
    assign proc_9_data_PIPO_blk[17] = 1'b0;
    assign proc_9_start_FIFO_blk[17] = 1'b0;
    assign proc_9_TLF_FIFO_blk[17] = 1'b0;
    assign proc_9_input_sync_blk[17] = 1'b0 | (ap_sync_load_value38_U0_ap_ready & load_value38_U0.ap_idle & ~ap_sync_load_value46_U0_ap_ready);
    assign proc_9_output_sync_blk[17] = 1'b0;
    assign proc_dep_vld_vec_9[17] = dl_detect_out ? proc_dep_vld_vec_9_reg[17] : (proc_9_data_FIFO_blk[17] | proc_9_data_PIPO_blk[17] | proc_9_start_FIFO_blk[17] | proc_9_TLF_FIFO_blk[17] | proc_9_input_sync_blk[17] | proc_9_output_sync_blk[17]);
    assign proc_9_data_FIFO_blk[18] = 1'b0;
    assign proc_9_data_PIPO_blk[18] = 1'b0;
    assign proc_9_start_FIFO_blk[18] = 1'b0;
    assign proc_9_TLF_FIFO_blk[18] = 1'b0;
    assign proc_9_input_sync_blk[18] = 1'b0 | (ap_sync_load_value38_U0_ap_ready & load_value38_U0.ap_idle & ~ap_sync_load_value47_U0_ap_ready);
    assign proc_9_output_sync_blk[18] = 1'b0;
    assign proc_dep_vld_vec_9[18] = dl_detect_out ? proc_dep_vld_vec_9_reg[18] : (proc_9_data_FIFO_blk[18] | proc_9_data_PIPO_blk[18] | proc_9_start_FIFO_blk[18] | proc_9_TLF_FIFO_blk[18] | proc_9_input_sync_blk[18] | proc_9_output_sync_blk[18]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_9_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_9_reg <= proc_dep_vld_vec_9;
        end
    end
    assign in_chan_dep_vld_vec_9[0] = dep_chan_vld_0_9;
    assign in_chan_dep_data_vec_9[34 : 0] = dep_chan_data_0_9;
    assign token_in_vec_9[0] = token_0_9;
    assign in_chan_dep_vld_vec_9[1] = dep_chan_vld_1_9;
    assign in_chan_dep_data_vec_9[69 : 35] = dep_chan_data_1_9;
    assign token_in_vec_9[1] = token_1_9;
    assign in_chan_dep_vld_vec_9[2] = dep_chan_vld_2_9;
    assign in_chan_dep_data_vec_9[104 : 70] = dep_chan_data_2_9;
    assign token_in_vec_9[2] = token_2_9;
    assign in_chan_dep_vld_vec_9[3] = dep_chan_vld_3_9;
    assign in_chan_dep_data_vec_9[139 : 105] = dep_chan_data_3_9;
    assign token_in_vec_9[3] = token_3_9;
    assign in_chan_dep_vld_vec_9[4] = dep_chan_vld_4_9;
    assign in_chan_dep_data_vec_9[174 : 140] = dep_chan_data_4_9;
    assign token_in_vec_9[4] = token_4_9;
    assign in_chan_dep_vld_vec_9[5] = dep_chan_vld_5_9;
    assign in_chan_dep_data_vec_9[209 : 175] = dep_chan_data_5_9;
    assign token_in_vec_9[5] = token_5_9;
    assign in_chan_dep_vld_vec_9[6] = dep_chan_vld_6_9;
    assign in_chan_dep_data_vec_9[244 : 210] = dep_chan_data_6_9;
    assign token_in_vec_9[6] = token_6_9;
    assign in_chan_dep_vld_vec_9[7] = dep_chan_vld_7_9;
    assign in_chan_dep_data_vec_9[279 : 245] = dep_chan_data_7_9;
    assign token_in_vec_9[7] = token_7_9;
    assign in_chan_dep_vld_vec_9[8] = dep_chan_vld_8_9;
    assign in_chan_dep_data_vec_9[314 : 280] = dep_chan_data_8_9;
    assign token_in_vec_9[8] = token_8_9;
    assign in_chan_dep_vld_vec_9[9] = dep_chan_vld_10_9;
    assign in_chan_dep_data_vec_9[349 : 315] = dep_chan_data_10_9;
    assign token_in_vec_9[9] = token_10_9;
    assign in_chan_dep_vld_vec_9[10] = dep_chan_vld_11_9;
    assign in_chan_dep_data_vec_9[384 : 350] = dep_chan_data_11_9;
    assign token_in_vec_9[10] = token_11_9;
    assign in_chan_dep_vld_vec_9[11] = dep_chan_vld_12_9;
    assign in_chan_dep_data_vec_9[419 : 385] = dep_chan_data_12_9;
    assign token_in_vec_9[11] = token_12_9;
    assign in_chan_dep_vld_vec_9[12] = dep_chan_vld_13_9;
    assign in_chan_dep_data_vec_9[454 : 420] = dep_chan_data_13_9;
    assign token_in_vec_9[12] = token_13_9;
    assign in_chan_dep_vld_vec_9[13] = dep_chan_vld_14_9;
    assign in_chan_dep_data_vec_9[489 : 455] = dep_chan_data_14_9;
    assign token_in_vec_9[13] = token_14_9;
    assign in_chan_dep_vld_vec_9[14] = dep_chan_vld_15_9;
    assign in_chan_dep_data_vec_9[524 : 490] = dep_chan_data_15_9;
    assign token_in_vec_9[14] = token_15_9;
    assign in_chan_dep_vld_vec_9[15] = dep_chan_vld_16_9;
    assign in_chan_dep_data_vec_9[559 : 525] = dep_chan_data_16_9;
    assign token_in_vec_9[15] = token_16_9;
    assign in_chan_dep_vld_vec_9[16] = dep_chan_vld_17_9;
    assign in_chan_dep_data_vec_9[594 : 560] = dep_chan_data_17_9;
    assign token_in_vec_9[16] = token_17_9;
    assign in_chan_dep_vld_vec_9[17] = dep_chan_vld_18_9;
    assign in_chan_dep_data_vec_9[629 : 595] = dep_chan_data_18_9;
    assign token_in_vec_9[17] = token_18_9;
    assign in_chan_dep_vld_vec_9[18] = dep_chan_vld_25_9;
    assign in_chan_dep_data_vec_9[664 : 630] = dep_chan_data_25_9;
    assign token_in_vec_9[18] = token_25_9;
    assign dep_chan_vld_9_0 = out_chan_dep_vld_vec_9[0];
    assign dep_chan_data_9_0 = out_chan_dep_data_9;
    assign token_9_0 = token_out_vec_9[0];
    assign dep_chan_vld_9_1 = out_chan_dep_vld_vec_9[1];
    assign dep_chan_data_9_1 = out_chan_dep_data_9;
    assign token_9_1 = token_out_vec_9[1];
    assign dep_chan_vld_9_25 = out_chan_dep_vld_vec_9[2];
    assign dep_chan_data_9_25 = out_chan_dep_data_9;
    assign token_9_25 = token_out_vec_9[2];
    assign dep_chan_vld_9_2 = out_chan_dep_vld_vec_9[3];
    assign dep_chan_data_9_2 = out_chan_dep_data_9;
    assign token_9_2 = token_out_vec_9[3];
    assign dep_chan_vld_9_3 = out_chan_dep_vld_vec_9[4];
    assign dep_chan_data_9_3 = out_chan_dep_data_9;
    assign token_9_3 = token_out_vec_9[4];
    assign dep_chan_vld_9_4 = out_chan_dep_vld_vec_9[5];
    assign dep_chan_data_9_4 = out_chan_dep_data_9;
    assign token_9_4 = token_out_vec_9[5];
    assign dep_chan_vld_9_5 = out_chan_dep_vld_vec_9[6];
    assign dep_chan_data_9_5 = out_chan_dep_data_9;
    assign token_9_5 = token_out_vec_9[6];
    assign dep_chan_vld_9_6 = out_chan_dep_vld_vec_9[7];
    assign dep_chan_data_9_6 = out_chan_dep_data_9;
    assign token_9_6 = token_out_vec_9[7];
    assign dep_chan_vld_9_7 = out_chan_dep_vld_vec_9[8];
    assign dep_chan_data_9_7 = out_chan_dep_data_9;
    assign token_9_7 = token_out_vec_9[8];
    assign dep_chan_vld_9_8 = out_chan_dep_vld_vec_9[9];
    assign dep_chan_data_9_8 = out_chan_dep_data_9;
    assign token_9_8 = token_out_vec_9[9];
    assign dep_chan_vld_9_10 = out_chan_dep_vld_vec_9[10];
    assign dep_chan_data_9_10 = out_chan_dep_data_9;
    assign token_9_10 = token_out_vec_9[10];
    assign dep_chan_vld_9_11 = out_chan_dep_vld_vec_9[11];
    assign dep_chan_data_9_11 = out_chan_dep_data_9;
    assign token_9_11 = token_out_vec_9[11];
    assign dep_chan_vld_9_12 = out_chan_dep_vld_vec_9[12];
    assign dep_chan_data_9_12 = out_chan_dep_data_9;
    assign token_9_12 = token_out_vec_9[12];
    assign dep_chan_vld_9_13 = out_chan_dep_vld_vec_9[13];
    assign dep_chan_data_9_13 = out_chan_dep_data_9;
    assign token_9_13 = token_out_vec_9[13];
    assign dep_chan_vld_9_14 = out_chan_dep_vld_vec_9[14];
    assign dep_chan_data_9_14 = out_chan_dep_data_9;
    assign token_9_14 = token_out_vec_9[14];
    assign dep_chan_vld_9_15 = out_chan_dep_vld_vec_9[15];
    assign dep_chan_data_9_15 = out_chan_dep_data_9;
    assign token_9_15 = token_out_vec_9[15];
    assign dep_chan_vld_9_16 = out_chan_dep_vld_vec_9[16];
    assign dep_chan_data_9_16 = out_chan_dep_data_9;
    assign token_9_16 = token_out_vec_9[16];
    assign dep_chan_vld_9_17 = out_chan_dep_vld_vec_9[17];
    assign dep_chan_data_9_17 = out_chan_dep_data_9;
    assign token_9_17 = token_out_vec_9[17];
    assign dep_chan_vld_9_18 = out_chan_dep_vld_vec_9[18];
    assign dep_chan_data_9_18 = out_chan_dep_data_9;
    assign token_9_18 = token_out_vec_9[18];

    // Process: load_value39_U0
    kernel_pr_hls_deadlock_detect_unit #(35, 10, 19, 19) kernel_pr_hls_deadlock_detect_unit_10 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_10),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_10),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_10),
        .token_in_vec(token_in_vec_10),
        .dl_detect_in(dl_detect_out),
        .origin(origin[10]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_10),
        .out_chan_dep_data(out_chan_dep_data_10),
        .token_out_vec(token_out_vec_10),
        .dl_detect_out(dl_in_vec[10]));

    assign proc_10_data_FIFO_blk[0] = 1'b0 | (~load_value39_U0.value_r_blk_n);
    assign proc_10_data_PIPO_blk[0] = 1'b0;
    assign proc_10_start_FIFO_blk[0] = 1'b0;
    assign proc_10_TLF_FIFO_blk[0] = 1'b0;
    assign proc_10_input_sync_blk[0] = 1'b0 | (ap_sync_load_value39_U0_ap_ready & load_value39_U0.ap_idle & ~ap_sync_kernel_pr_entry98_U0_ap_ready);
    assign proc_10_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_10[0] = dl_detect_out ? proc_dep_vld_vec_10_reg[0] : (proc_10_data_FIFO_blk[0] | proc_10_data_PIPO_blk[0] | proc_10_start_FIFO_blk[0] | proc_10_TLF_FIFO_blk[0] | proc_10_input_sync_blk[0] | proc_10_output_sync_blk[0]);
    assign proc_10_data_FIFO_blk[1] = 1'b0 | (~load_value39_U0.bipedge_size_blk_n) | (~load_value39_U0.bipedge_stream_V_V7_blk_n);
    assign proc_10_data_PIPO_blk[1] = 1'b0;
    assign proc_10_start_FIFO_blk[1] = 1'b0;
    assign proc_10_TLF_FIFO_blk[1] = 1'b0;
    assign proc_10_input_sync_blk[1] = 1'b0 | (ap_sync_load_value39_U0_ap_ready & load_value39_U0.ap_idle & ~ap_sync_load_bipedge30_U0_ap_ready);
    assign proc_10_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_10[1] = dl_detect_out ? proc_dep_vld_vec_10_reg[1] : (proc_10_data_FIFO_blk[1] | proc_10_data_PIPO_blk[1] | proc_10_start_FIFO_blk[1] | proc_10_TLF_FIFO_blk[1] | proc_10_input_sync_blk[1] | proc_10_output_sync_blk[1]);
    assign proc_10_data_FIFO_blk[2] = 1'b0 | (~load_value39_U0.value_stream_V_V22_blk_n);
    assign proc_10_data_PIPO_blk[2] = 1'b0;
    assign proc_10_start_FIFO_blk[2] = 1'b0;
    assign proc_10_TLF_FIFO_blk[2] = 1'b0;
    assign proc_10_input_sync_blk[2] = 1'b0;
    assign proc_10_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_10[2] = dl_detect_out ? proc_dep_vld_vec_10_reg[2] : (proc_10_data_FIFO_blk[2] | proc_10_data_PIPO_blk[2] | proc_10_start_FIFO_blk[2] | proc_10_TLF_FIFO_blk[2] | proc_10_input_sync_blk[2] | proc_10_output_sync_blk[2]);
    assign proc_10_data_FIFO_blk[3] = 1'b0;
    assign proc_10_data_PIPO_blk[3] = 1'b0;
    assign proc_10_start_FIFO_blk[3] = 1'b0;
    assign proc_10_TLF_FIFO_blk[3] = 1'b0;
    assign proc_10_input_sync_blk[3] = 1'b0 | (ap_sync_load_value39_U0_ap_ready & load_value39_U0.ap_idle & ~ap_sync_load_bipedge31_U0_ap_ready);
    assign proc_10_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_10[3] = dl_detect_out ? proc_dep_vld_vec_10_reg[3] : (proc_10_data_FIFO_blk[3] | proc_10_data_PIPO_blk[3] | proc_10_start_FIFO_blk[3] | proc_10_TLF_FIFO_blk[3] | proc_10_input_sync_blk[3] | proc_10_output_sync_blk[3]);
    assign proc_10_data_FIFO_blk[4] = 1'b0;
    assign proc_10_data_PIPO_blk[4] = 1'b0;
    assign proc_10_start_FIFO_blk[4] = 1'b0;
    assign proc_10_TLF_FIFO_blk[4] = 1'b0;
    assign proc_10_input_sync_blk[4] = 1'b0 | (ap_sync_load_value39_U0_ap_ready & load_value39_U0.ap_idle & ~ap_sync_load_value32_U0_ap_ready);
    assign proc_10_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_10[4] = dl_detect_out ? proc_dep_vld_vec_10_reg[4] : (proc_10_data_FIFO_blk[4] | proc_10_data_PIPO_blk[4] | proc_10_start_FIFO_blk[4] | proc_10_TLF_FIFO_blk[4] | proc_10_input_sync_blk[4] | proc_10_output_sync_blk[4]);
    assign proc_10_data_FIFO_blk[5] = 1'b0;
    assign proc_10_data_PIPO_blk[5] = 1'b0;
    assign proc_10_start_FIFO_blk[5] = 1'b0;
    assign proc_10_TLF_FIFO_blk[5] = 1'b0;
    assign proc_10_input_sync_blk[5] = 1'b0 | (ap_sync_load_value39_U0_ap_ready & load_value39_U0.ap_idle & ~ap_sync_load_value33_U0_ap_ready);
    assign proc_10_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_10[5] = dl_detect_out ? proc_dep_vld_vec_10_reg[5] : (proc_10_data_FIFO_blk[5] | proc_10_data_PIPO_blk[5] | proc_10_start_FIFO_blk[5] | proc_10_TLF_FIFO_blk[5] | proc_10_input_sync_blk[5] | proc_10_output_sync_blk[5]);
    assign proc_10_data_FIFO_blk[6] = 1'b0;
    assign proc_10_data_PIPO_blk[6] = 1'b0;
    assign proc_10_start_FIFO_blk[6] = 1'b0;
    assign proc_10_TLF_FIFO_blk[6] = 1'b0;
    assign proc_10_input_sync_blk[6] = 1'b0 | (ap_sync_load_value39_U0_ap_ready & load_value39_U0.ap_idle & ~ap_sync_load_value34_U0_ap_ready);
    assign proc_10_output_sync_blk[6] = 1'b0;
    assign proc_dep_vld_vec_10[6] = dl_detect_out ? proc_dep_vld_vec_10_reg[6] : (proc_10_data_FIFO_blk[6] | proc_10_data_PIPO_blk[6] | proc_10_start_FIFO_blk[6] | proc_10_TLF_FIFO_blk[6] | proc_10_input_sync_blk[6] | proc_10_output_sync_blk[6]);
    assign proc_10_data_FIFO_blk[7] = 1'b0;
    assign proc_10_data_PIPO_blk[7] = 1'b0;
    assign proc_10_start_FIFO_blk[7] = 1'b0;
    assign proc_10_TLF_FIFO_blk[7] = 1'b0;
    assign proc_10_input_sync_blk[7] = 1'b0 | (ap_sync_load_value39_U0_ap_ready & load_value39_U0.ap_idle & ~ap_sync_load_value35_U0_ap_ready);
    assign proc_10_output_sync_blk[7] = 1'b0;
    assign proc_dep_vld_vec_10[7] = dl_detect_out ? proc_dep_vld_vec_10_reg[7] : (proc_10_data_FIFO_blk[7] | proc_10_data_PIPO_blk[7] | proc_10_start_FIFO_blk[7] | proc_10_TLF_FIFO_blk[7] | proc_10_input_sync_blk[7] | proc_10_output_sync_blk[7]);
    assign proc_10_data_FIFO_blk[8] = 1'b0;
    assign proc_10_data_PIPO_blk[8] = 1'b0;
    assign proc_10_start_FIFO_blk[8] = 1'b0;
    assign proc_10_TLF_FIFO_blk[8] = 1'b0;
    assign proc_10_input_sync_blk[8] = 1'b0 | (ap_sync_load_value39_U0_ap_ready & load_value39_U0.ap_idle & ~ap_sync_load_value36_U0_ap_ready);
    assign proc_10_output_sync_blk[8] = 1'b0;
    assign proc_dep_vld_vec_10[8] = dl_detect_out ? proc_dep_vld_vec_10_reg[8] : (proc_10_data_FIFO_blk[8] | proc_10_data_PIPO_blk[8] | proc_10_start_FIFO_blk[8] | proc_10_TLF_FIFO_blk[8] | proc_10_input_sync_blk[8] | proc_10_output_sync_blk[8]);
    assign proc_10_data_FIFO_blk[9] = 1'b0;
    assign proc_10_data_PIPO_blk[9] = 1'b0;
    assign proc_10_start_FIFO_blk[9] = 1'b0;
    assign proc_10_TLF_FIFO_blk[9] = 1'b0;
    assign proc_10_input_sync_blk[9] = 1'b0 | (ap_sync_load_value39_U0_ap_ready & load_value39_U0.ap_idle & ~ap_sync_load_value37_U0_ap_ready);
    assign proc_10_output_sync_blk[9] = 1'b0;
    assign proc_dep_vld_vec_10[9] = dl_detect_out ? proc_dep_vld_vec_10_reg[9] : (proc_10_data_FIFO_blk[9] | proc_10_data_PIPO_blk[9] | proc_10_start_FIFO_blk[9] | proc_10_TLF_FIFO_blk[9] | proc_10_input_sync_blk[9] | proc_10_output_sync_blk[9]);
    assign proc_10_data_FIFO_blk[10] = 1'b0;
    assign proc_10_data_PIPO_blk[10] = 1'b0;
    assign proc_10_start_FIFO_blk[10] = 1'b0;
    assign proc_10_TLF_FIFO_blk[10] = 1'b0;
    assign proc_10_input_sync_blk[10] = 1'b0 | (ap_sync_load_value39_U0_ap_ready & load_value39_U0.ap_idle & ~ap_sync_load_value38_U0_ap_ready);
    assign proc_10_output_sync_blk[10] = 1'b0;
    assign proc_dep_vld_vec_10[10] = dl_detect_out ? proc_dep_vld_vec_10_reg[10] : (proc_10_data_FIFO_blk[10] | proc_10_data_PIPO_blk[10] | proc_10_start_FIFO_blk[10] | proc_10_TLF_FIFO_blk[10] | proc_10_input_sync_blk[10] | proc_10_output_sync_blk[10]);
    assign proc_10_data_FIFO_blk[11] = 1'b0;
    assign proc_10_data_PIPO_blk[11] = 1'b0;
    assign proc_10_start_FIFO_blk[11] = 1'b0;
    assign proc_10_TLF_FIFO_blk[11] = 1'b0;
    assign proc_10_input_sync_blk[11] = 1'b0 | (ap_sync_load_value39_U0_ap_ready & load_value39_U0.ap_idle & ~ap_sync_load_value40_U0_ap_ready);
    assign proc_10_output_sync_blk[11] = 1'b0;
    assign proc_dep_vld_vec_10[11] = dl_detect_out ? proc_dep_vld_vec_10_reg[11] : (proc_10_data_FIFO_blk[11] | proc_10_data_PIPO_blk[11] | proc_10_start_FIFO_blk[11] | proc_10_TLF_FIFO_blk[11] | proc_10_input_sync_blk[11] | proc_10_output_sync_blk[11]);
    assign proc_10_data_FIFO_blk[12] = 1'b0;
    assign proc_10_data_PIPO_blk[12] = 1'b0;
    assign proc_10_start_FIFO_blk[12] = 1'b0;
    assign proc_10_TLF_FIFO_blk[12] = 1'b0;
    assign proc_10_input_sync_blk[12] = 1'b0 | (ap_sync_load_value39_U0_ap_ready & load_value39_U0.ap_idle & ~ap_sync_load_value41_U0_ap_ready);
    assign proc_10_output_sync_blk[12] = 1'b0;
    assign proc_dep_vld_vec_10[12] = dl_detect_out ? proc_dep_vld_vec_10_reg[12] : (proc_10_data_FIFO_blk[12] | proc_10_data_PIPO_blk[12] | proc_10_start_FIFO_blk[12] | proc_10_TLF_FIFO_blk[12] | proc_10_input_sync_blk[12] | proc_10_output_sync_blk[12]);
    assign proc_10_data_FIFO_blk[13] = 1'b0;
    assign proc_10_data_PIPO_blk[13] = 1'b0;
    assign proc_10_start_FIFO_blk[13] = 1'b0;
    assign proc_10_TLF_FIFO_blk[13] = 1'b0;
    assign proc_10_input_sync_blk[13] = 1'b0 | (ap_sync_load_value39_U0_ap_ready & load_value39_U0.ap_idle & ~ap_sync_load_value42_U0_ap_ready);
    assign proc_10_output_sync_blk[13] = 1'b0;
    assign proc_dep_vld_vec_10[13] = dl_detect_out ? proc_dep_vld_vec_10_reg[13] : (proc_10_data_FIFO_blk[13] | proc_10_data_PIPO_blk[13] | proc_10_start_FIFO_blk[13] | proc_10_TLF_FIFO_blk[13] | proc_10_input_sync_blk[13] | proc_10_output_sync_blk[13]);
    assign proc_10_data_FIFO_blk[14] = 1'b0;
    assign proc_10_data_PIPO_blk[14] = 1'b0;
    assign proc_10_start_FIFO_blk[14] = 1'b0;
    assign proc_10_TLF_FIFO_blk[14] = 1'b0;
    assign proc_10_input_sync_blk[14] = 1'b0 | (ap_sync_load_value39_U0_ap_ready & load_value39_U0.ap_idle & ~ap_sync_load_value43_U0_ap_ready);
    assign proc_10_output_sync_blk[14] = 1'b0;
    assign proc_dep_vld_vec_10[14] = dl_detect_out ? proc_dep_vld_vec_10_reg[14] : (proc_10_data_FIFO_blk[14] | proc_10_data_PIPO_blk[14] | proc_10_start_FIFO_blk[14] | proc_10_TLF_FIFO_blk[14] | proc_10_input_sync_blk[14] | proc_10_output_sync_blk[14]);
    assign proc_10_data_FIFO_blk[15] = 1'b0;
    assign proc_10_data_PIPO_blk[15] = 1'b0;
    assign proc_10_start_FIFO_blk[15] = 1'b0;
    assign proc_10_TLF_FIFO_blk[15] = 1'b0;
    assign proc_10_input_sync_blk[15] = 1'b0 | (ap_sync_load_value39_U0_ap_ready & load_value39_U0.ap_idle & ~ap_sync_load_value44_U0_ap_ready);
    assign proc_10_output_sync_blk[15] = 1'b0;
    assign proc_dep_vld_vec_10[15] = dl_detect_out ? proc_dep_vld_vec_10_reg[15] : (proc_10_data_FIFO_blk[15] | proc_10_data_PIPO_blk[15] | proc_10_start_FIFO_blk[15] | proc_10_TLF_FIFO_blk[15] | proc_10_input_sync_blk[15] | proc_10_output_sync_blk[15]);
    assign proc_10_data_FIFO_blk[16] = 1'b0;
    assign proc_10_data_PIPO_blk[16] = 1'b0;
    assign proc_10_start_FIFO_blk[16] = 1'b0;
    assign proc_10_TLF_FIFO_blk[16] = 1'b0;
    assign proc_10_input_sync_blk[16] = 1'b0 | (ap_sync_load_value39_U0_ap_ready & load_value39_U0.ap_idle & ~ap_sync_load_value45_U0_ap_ready);
    assign proc_10_output_sync_blk[16] = 1'b0;
    assign proc_dep_vld_vec_10[16] = dl_detect_out ? proc_dep_vld_vec_10_reg[16] : (proc_10_data_FIFO_blk[16] | proc_10_data_PIPO_blk[16] | proc_10_start_FIFO_blk[16] | proc_10_TLF_FIFO_blk[16] | proc_10_input_sync_blk[16] | proc_10_output_sync_blk[16]);
    assign proc_10_data_FIFO_blk[17] = 1'b0;
    assign proc_10_data_PIPO_blk[17] = 1'b0;
    assign proc_10_start_FIFO_blk[17] = 1'b0;
    assign proc_10_TLF_FIFO_blk[17] = 1'b0;
    assign proc_10_input_sync_blk[17] = 1'b0 | (ap_sync_load_value39_U0_ap_ready & load_value39_U0.ap_idle & ~ap_sync_load_value46_U0_ap_ready);
    assign proc_10_output_sync_blk[17] = 1'b0;
    assign proc_dep_vld_vec_10[17] = dl_detect_out ? proc_dep_vld_vec_10_reg[17] : (proc_10_data_FIFO_blk[17] | proc_10_data_PIPO_blk[17] | proc_10_start_FIFO_blk[17] | proc_10_TLF_FIFO_blk[17] | proc_10_input_sync_blk[17] | proc_10_output_sync_blk[17]);
    assign proc_10_data_FIFO_blk[18] = 1'b0;
    assign proc_10_data_PIPO_blk[18] = 1'b0;
    assign proc_10_start_FIFO_blk[18] = 1'b0;
    assign proc_10_TLF_FIFO_blk[18] = 1'b0;
    assign proc_10_input_sync_blk[18] = 1'b0 | (ap_sync_load_value39_U0_ap_ready & load_value39_U0.ap_idle & ~ap_sync_load_value47_U0_ap_ready);
    assign proc_10_output_sync_blk[18] = 1'b0;
    assign proc_dep_vld_vec_10[18] = dl_detect_out ? proc_dep_vld_vec_10_reg[18] : (proc_10_data_FIFO_blk[18] | proc_10_data_PIPO_blk[18] | proc_10_start_FIFO_blk[18] | proc_10_TLF_FIFO_blk[18] | proc_10_input_sync_blk[18] | proc_10_output_sync_blk[18]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_10_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_10_reg <= proc_dep_vld_vec_10;
        end
    end
    assign in_chan_dep_vld_vec_10[0] = dep_chan_vld_0_10;
    assign in_chan_dep_data_vec_10[34 : 0] = dep_chan_data_0_10;
    assign token_in_vec_10[0] = token_0_10;
    assign in_chan_dep_vld_vec_10[1] = dep_chan_vld_1_10;
    assign in_chan_dep_data_vec_10[69 : 35] = dep_chan_data_1_10;
    assign token_in_vec_10[1] = token_1_10;
    assign in_chan_dep_vld_vec_10[2] = dep_chan_vld_2_10;
    assign in_chan_dep_data_vec_10[104 : 70] = dep_chan_data_2_10;
    assign token_in_vec_10[2] = token_2_10;
    assign in_chan_dep_vld_vec_10[3] = dep_chan_vld_3_10;
    assign in_chan_dep_data_vec_10[139 : 105] = dep_chan_data_3_10;
    assign token_in_vec_10[3] = token_3_10;
    assign in_chan_dep_vld_vec_10[4] = dep_chan_vld_4_10;
    assign in_chan_dep_data_vec_10[174 : 140] = dep_chan_data_4_10;
    assign token_in_vec_10[4] = token_4_10;
    assign in_chan_dep_vld_vec_10[5] = dep_chan_vld_5_10;
    assign in_chan_dep_data_vec_10[209 : 175] = dep_chan_data_5_10;
    assign token_in_vec_10[5] = token_5_10;
    assign in_chan_dep_vld_vec_10[6] = dep_chan_vld_6_10;
    assign in_chan_dep_data_vec_10[244 : 210] = dep_chan_data_6_10;
    assign token_in_vec_10[6] = token_6_10;
    assign in_chan_dep_vld_vec_10[7] = dep_chan_vld_7_10;
    assign in_chan_dep_data_vec_10[279 : 245] = dep_chan_data_7_10;
    assign token_in_vec_10[7] = token_7_10;
    assign in_chan_dep_vld_vec_10[8] = dep_chan_vld_8_10;
    assign in_chan_dep_data_vec_10[314 : 280] = dep_chan_data_8_10;
    assign token_in_vec_10[8] = token_8_10;
    assign in_chan_dep_vld_vec_10[9] = dep_chan_vld_9_10;
    assign in_chan_dep_data_vec_10[349 : 315] = dep_chan_data_9_10;
    assign token_in_vec_10[9] = token_9_10;
    assign in_chan_dep_vld_vec_10[10] = dep_chan_vld_11_10;
    assign in_chan_dep_data_vec_10[384 : 350] = dep_chan_data_11_10;
    assign token_in_vec_10[10] = token_11_10;
    assign in_chan_dep_vld_vec_10[11] = dep_chan_vld_12_10;
    assign in_chan_dep_data_vec_10[419 : 385] = dep_chan_data_12_10;
    assign token_in_vec_10[11] = token_12_10;
    assign in_chan_dep_vld_vec_10[12] = dep_chan_vld_13_10;
    assign in_chan_dep_data_vec_10[454 : 420] = dep_chan_data_13_10;
    assign token_in_vec_10[12] = token_13_10;
    assign in_chan_dep_vld_vec_10[13] = dep_chan_vld_14_10;
    assign in_chan_dep_data_vec_10[489 : 455] = dep_chan_data_14_10;
    assign token_in_vec_10[13] = token_14_10;
    assign in_chan_dep_vld_vec_10[14] = dep_chan_vld_15_10;
    assign in_chan_dep_data_vec_10[524 : 490] = dep_chan_data_15_10;
    assign token_in_vec_10[14] = token_15_10;
    assign in_chan_dep_vld_vec_10[15] = dep_chan_vld_16_10;
    assign in_chan_dep_data_vec_10[559 : 525] = dep_chan_data_16_10;
    assign token_in_vec_10[15] = token_16_10;
    assign in_chan_dep_vld_vec_10[16] = dep_chan_vld_17_10;
    assign in_chan_dep_data_vec_10[594 : 560] = dep_chan_data_17_10;
    assign token_in_vec_10[16] = token_17_10;
    assign in_chan_dep_vld_vec_10[17] = dep_chan_vld_18_10;
    assign in_chan_dep_data_vec_10[629 : 595] = dep_chan_data_18_10;
    assign token_in_vec_10[17] = token_18_10;
    assign in_chan_dep_vld_vec_10[18] = dep_chan_vld_26_10;
    assign in_chan_dep_data_vec_10[664 : 630] = dep_chan_data_26_10;
    assign token_in_vec_10[18] = token_26_10;
    assign dep_chan_vld_10_0 = out_chan_dep_vld_vec_10[0];
    assign dep_chan_data_10_0 = out_chan_dep_data_10;
    assign token_10_0 = token_out_vec_10[0];
    assign dep_chan_vld_10_1 = out_chan_dep_vld_vec_10[1];
    assign dep_chan_data_10_1 = out_chan_dep_data_10;
    assign token_10_1 = token_out_vec_10[1];
    assign dep_chan_vld_10_26 = out_chan_dep_vld_vec_10[2];
    assign dep_chan_data_10_26 = out_chan_dep_data_10;
    assign token_10_26 = token_out_vec_10[2];
    assign dep_chan_vld_10_2 = out_chan_dep_vld_vec_10[3];
    assign dep_chan_data_10_2 = out_chan_dep_data_10;
    assign token_10_2 = token_out_vec_10[3];
    assign dep_chan_vld_10_3 = out_chan_dep_vld_vec_10[4];
    assign dep_chan_data_10_3 = out_chan_dep_data_10;
    assign token_10_3 = token_out_vec_10[4];
    assign dep_chan_vld_10_4 = out_chan_dep_vld_vec_10[5];
    assign dep_chan_data_10_4 = out_chan_dep_data_10;
    assign token_10_4 = token_out_vec_10[5];
    assign dep_chan_vld_10_5 = out_chan_dep_vld_vec_10[6];
    assign dep_chan_data_10_5 = out_chan_dep_data_10;
    assign token_10_5 = token_out_vec_10[6];
    assign dep_chan_vld_10_6 = out_chan_dep_vld_vec_10[7];
    assign dep_chan_data_10_6 = out_chan_dep_data_10;
    assign token_10_6 = token_out_vec_10[7];
    assign dep_chan_vld_10_7 = out_chan_dep_vld_vec_10[8];
    assign dep_chan_data_10_7 = out_chan_dep_data_10;
    assign token_10_7 = token_out_vec_10[8];
    assign dep_chan_vld_10_8 = out_chan_dep_vld_vec_10[9];
    assign dep_chan_data_10_8 = out_chan_dep_data_10;
    assign token_10_8 = token_out_vec_10[9];
    assign dep_chan_vld_10_9 = out_chan_dep_vld_vec_10[10];
    assign dep_chan_data_10_9 = out_chan_dep_data_10;
    assign token_10_9 = token_out_vec_10[10];
    assign dep_chan_vld_10_11 = out_chan_dep_vld_vec_10[11];
    assign dep_chan_data_10_11 = out_chan_dep_data_10;
    assign token_10_11 = token_out_vec_10[11];
    assign dep_chan_vld_10_12 = out_chan_dep_vld_vec_10[12];
    assign dep_chan_data_10_12 = out_chan_dep_data_10;
    assign token_10_12 = token_out_vec_10[12];
    assign dep_chan_vld_10_13 = out_chan_dep_vld_vec_10[13];
    assign dep_chan_data_10_13 = out_chan_dep_data_10;
    assign token_10_13 = token_out_vec_10[13];
    assign dep_chan_vld_10_14 = out_chan_dep_vld_vec_10[14];
    assign dep_chan_data_10_14 = out_chan_dep_data_10;
    assign token_10_14 = token_out_vec_10[14];
    assign dep_chan_vld_10_15 = out_chan_dep_vld_vec_10[15];
    assign dep_chan_data_10_15 = out_chan_dep_data_10;
    assign token_10_15 = token_out_vec_10[15];
    assign dep_chan_vld_10_16 = out_chan_dep_vld_vec_10[16];
    assign dep_chan_data_10_16 = out_chan_dep_data_10;
    assign token_10_16 = token_out_vec_10[16];
    assign dep_chan_vld_10_17 = out_chan_dep_vld_vec_10[17];
    assign dep_chan_data_10_17 = out_chan_dep_data_10;
    assign token_10_17 = token_out_vec_10[17];
    assign dep_chan_vld_10_18 = out_chan_dep_vld_vec_10[18];
    assign dep_chan_data_10_18 = out_chan_dep_data_10;
    assign token_10_18 = token_out_vec_10[18];

    // Process: load_value40_U0
    kernel_pr_hls_deadlock_detect_unit #(35, 11, 19, 19) kernel_pr_hls_deadlock_detect_unit_11 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_11),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_11),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_11),
        .token_in_vec(token_in_vec_11),
        .dl_detect_in(dl_detect_out),
        .origin(origin[11]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_11),
        .out_chan_dep_data(out_chan_dep_data_11),
        .token_out_vec(token_out_vec_11),
        .dl_detect_out(dl_in_vec[11]));

    assign proc_11_data_FIFO_blk[0] = 1'b0 | (~load_value40_U0.value_r_blk_n);
    assign proc_11_data_PIPO_blk[0] = 1'b0;
    assign proc_11_start_FIFO_blk[0] = 1'b0;
    assign proc_11_TLF_FIFO_blk[0] = 1'b0;
    assign proc_11_input_sync_blk[0] = 1'b0 | (ap_sync_load_value40_U0_ap_ready & load_value40_U0.ap_idle & ~ap_sync_kernel_pr_entry98_U0_ap_ready);
    assign proc_11_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_11[0] = dl_detect_out ? proc_dep_vld_vec_11_reg[0] : (proc_11_data_FIFO_blk[0] | proc_11_data_PIPO_blk[0] | proc_11_start_FIFO_blk[0] | proc_11_TLF_FIFO_blk[0] | proc_11_input_sync_blk[0] | proc_11_output_sync_blk[0]);
    assign proc_11_data_FIFO_blk[1] = 1'b0 | (~load_value40_U0.bipedge_size_blk_n) | (~load_value40_U0.bipedge_stream_V_V8_blk_n);
    assign proc_11_data_PIPO_blk[1] = 1'b0;
    assign proc_11_start_FIFO_blk[1] = 1'b0;
    assign proc_11_TLF_FIFO_blk[1] = 1'b0;
    assign proc_11_input_sync_blk[1] = 1'b0 | (ap_sync_load_value40_U0_ap_ready & load_value40_U0.ap_idle & ~ap_sync_load_bipedge31_U0_ap_ready);
    assign proc_11_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_11[1] = dl_detect_out ? proc_dep_vld_vec_11_reg[1] : (proc_11_data_FIFO_blk[1] | proc_11_data_PIPO_blk[1] | proc_11_start_FIFO_blk[1] | proc_11_TLF_FIFO_blk[1] | proc_11_input_sync_blk[1] | proc_11_output_sync_blk[1]);
    assign proc_11_data_FIFO_blk[2] = 1'b0 | (~load_value40_U0.value_stream_V_V23_blk_n);
    assign proc_11_data_PIPO_blk[2] = 1'b0;
    assign proc_11_start_FIFO_blk[2] = 1'b0;
    assign proc_11_TLF_FIFO_blk[2] = 1'b0;
    assign proc_11_input_sync_blk[2] = 1'b0;
    assign proc_11_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_11[2] = dl_detect_out ? proc_dep_vld_vec_11_reg[2] : (proc_11_data_FIFO_blk[2] | proc_11_data_PIPO_blk[2] | proc_11_start_FIFO_blk[2] | proc_11_TLF_FIFO_blk[2] | proc_11_input_sync_blk[2] | proc_11_output_sync_blk[2]);
    assign proc_11_data_FIFO_blk[3] = 1'b0;
    assign proc_11_data_PIPO_blk[3] = 1'b0;
    assign proc_11_start_FIFO_blk[3] = 1'b0;
    assign proc_11_TLF_FIFO_blk[3] = 1'b0;
    assign proc_11_input_sync_blk[3] = 1'b0 | (ap_sync_load_value40_U0_ap_ready & load_value40_U0.ap_idle & ~ap_sync_load_bipedge30_U0_ap_ready);
    assign proc_11_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_11[3] = dl_detect_out ? proc_dep_vld_vec_11_reg[3] : (proc_11_data_FIFO_blk[3] | proc_11_data_PIPO_blk[3] | proc_11_start_FIFO_blk[3] | proc_11_TLF_FIFO_blk[3] | proc_11_input_sync_blk[3] | proc_11_output_sync_blk[3]);
    assign proc_11_data_FIFO_blk[4] = 1'b0;
    assign proc_11_data_PIPO_blk[4] = 1'b0;
    assign proc_11_start_FIFO_blk[4] = 1'b0;
    assign proc_11_TLF_FIFO_blk[4] = 1'b0;
    assign proc_11_input_sync_blk[4] = 1'b0 | (ap_sync_load_value40_U0_ap_ready & load_value40_U0.ap_idle & ~ap_sync_load_value32_U0_ap_ready);
    assign proc_11_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_11[4] = dl_detect_out ? proc_dep_vld_vec_11_reg[4] : (proc_11_data_FIFO_blk[4] | proc_11_data_PIPO_blk[4] | proc_11_start_FIFO_blk[4] | proc_11_TLF_FIFO_blk[4] | proc_11_input_sync_blk[4] | proc_11_output_sync_blk[4]);
    assign proc_11_data_FIFO_blk[5] = 1'b0;
    assign proc_11_data_PIPO_blk[5] = 1'b0;
    assign proc_11_start_FIFO_blk[5] = 1'b0;
    assign proc_11_TLF_FIFO_blk[5] = 1'b0;
    assign proc_11_input_sync_blk[5] = 1'b0 | (ap_sync_load_value40_U0_ap_ready & load_value40_U0.ap_idle & ~ap_sync_load_value33_U0_ap_ready);
    assign proc_11_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_11[5] = dl_detect_out ? proc_dep_vld_vec_11_reg[5] : (proc_11_data_FIFO_blk[5] | proc_11_data_PIPO_blk[5] | proc_11_start_FIFO_blk[5] | proc_11_TLF_FIFO_blk[5] | proc_11_input_sync_blk[5] | proc_11_output_sync_blk[5]);
    assign proc_11_data_FIFO_blk[6] = 1'b0;
    assign proc_11_data_PIPO_blk[6] = 1'b0;
    assign proc_11_start_FIFO_blk[6] = 1'b0;
    assign proc_11_TLF_FIFO_blk[6] = 1'b0;
    assign proc_11_input_sync_blk[6] = 1'b0 | (ap_sync_load_value40_U0_ap_ready & load_value40_U0.ap_idle & ~ap_sync_load_value34_U0_ap_ready);
    assign proc_11_output_sync_blk[6] = 1'b0;
    assign proc_dep_vld_vec_11[6] = dl_detect_out ? proc_dep_vld_vec_11_reg[6] : (proc_11_data_FIFO_blk[6] | proc_11_data_PIPO_blk[6] | proc_11_start_FIFO_blk[6] | proc_11_TLF_FIFO_blk[6] | proc_11_input_sync_blk[6] | proc_11_output_sync_blk[6]);
    assign proc_11_data_FIFO_blk[7] = 1'b0;
    assign proc_11_data_PIPO_blk[7] = 1'b0;
    assign proc_11_start_FIFO_blk[7] = 1'b0;
    assign proc_11_TLF_FIFO_blk[7] = 1'b0;
    assign proc_11_input_sync_blk[7] = 1'b0 | (ap_sync_load_value40_U0_ap_ready & load_value40_U0.ap_idle & ~ap_sync_load_value35_U0_ap_ready);
    assign proc_11_output_sync_blk[7] = 1'b0;
    assign proc_dep_vld_vec_11[7] = dl_detect_out ? proc_dep_vld_vec_11_reg[7] : (proc_11_data_FIFO_blk[7] | proc_11_data_PIPO_blk[7] | proc_11_start_FIFO_blk[7] | proc_11_TLF_FIFO_blk[7] | proc_11_input_sync_blk[7] | proc_11_output_sync_blk[7]);
    assign proc_11_data_FIFO_blk[8] = 1'b0;
    assign proc_11_data_PIPO_blk[8] = 1'b0;
    assign proc_11_start_FIFO_blk[8] = 1'b0;
    assign proc_11_TLF_FIFO_blk[8] = 1'b0;
    assign proc_11_input_sync_blk[8] = 1'b0 | (ap_sync_load_value40_U0_ap_ready & load_value40_U0.ap_idle & ~ap_sync_load_value36_U0_ap_ready);
    assign proc_11_output_sync_blk[8] = 1'b0;
    assign proc_dep_vld_vec_11[8] = dl_detect_out ? proc_dep_vld_vec_11_reg[8] : (proc_11_data_FIFO_blk[8] | proc_11_data_PIPO_blk[8] | proc_11_start_FIFO_blk[8] | proc_11_TLF_FIFO_blk[8] | proc_11_input_sync_blk[8] | proc_11_output_sync_blk[8]);
    assign proc_11_data_FIFO_blk[9] = 1'b0;
    assign proc_11_data_PIPO_blk[9] = 1'b0;
    assign proc_11_start_FIFO_blk[9] = 1'b0;
    assign proc_11_TLF_FIFO_blk[9] = 1'b0;
    assign proc_11_input_sync_blk[9] = 1'b0 | (ap_sync_load_value40_U0_ap_ready & load_value40_U0.ap_idle & ~ap_sync_load_value37_U0_ap_ready);
    assign proc_11_output_sync_blk[9] = 1'b0;
    assign proc_dep_vld_vec_11[9] = dl_detect_out ? proc_dep_vld_vec_11_reg[9] : (proc_11_data_FIFO_blk[9] | proc_11_data_PIPO_blk[9] | proc_11_start_FIFO_blk[9] | proc_11_TLF_FIFO_blk[9] | proc_11_input_sync_blk[9] | proc_11_output_sync_blk[9]);
    assign proc_11_data_FIFO_blk[10] = 1'b0;
    assign proc_11_data_PIPO_blk[10] = 1'b0;
    assign proc_11_start_FIFO_blk[10] = 1'b0;
    assign proc_11_TLF_FIFO_blk[10] = 1'b0;
    assign proc_11_input_sync_blk[10] = 1'b0 | (ap_sync_load_value40_U0_ap_ready & load_value40_U0.ap_idle & ~ap_sync_load_value38_U0_ap_ready);
    assign proc_11_output_sync_blk[10] = 1'b0;
    assign proc_dep_vld_vec_11[10] = dl_detect_out ? proc_dep_vld_vec_11_reg[10] : (proc_11_data_FIFO_blk[10] | proc_11_data_PIPO_blk[10] | proc_11_start_FIFO_blk[10] | proc_11_TLF_FIFO_blk[10] | proc_11_input_sync_blk[10] | proc_11_output_sync_blk[10]);
    assign proc_11_data_FIFO_blk[11] = 1'b0;
    assign proc_11_data_PIPO_blk[11] = 1'b0;
    assign proc_11_start_FIFO_blk[11] = 1'b0;
    assign proc_11_TLF_FIFO_blk[11] = 1'b0;
    assign proc_11_input_sync_blk[11] = 1'b0 | (ap_sync_load_value40_U0_ap_ready & load_value40_U0.ap_idle & ~ap_sync_load_value39_U0_ap_ready);
    assign proc_11_output_sync_blk[11] = 1'b0;
    assign proc_dep_vld_vec_11[11] = dl_detect_out ? proc_dep_vld_vec_11_reg[11] : (proc_11_data_FIFO_blk[11] | proc_11_data_PIPO_blk[11] | proc_11_start_FIFO_blk[11] | proc_11_TLF_FIFO_blk[11] | proc_11_input_sync_blk[11] | proc_11_output_sync_blk[11]);
    assign proc_11_data_FIFO_blk[12] = 1'b0;
    assign proc_11_data_PIPO_blk[12] = 1'b0;
    assign proc_11_start_FIFO_blk[12] = 1'b0;
    assign proc_11_TLF_FIFO_blk[12] = 1'b0;
    assign proc_11_input_sync_blk[12] = 1'b0 | (ap_sync_load_value40_U0_ap_ready & load_value40_U0.ap_idle & ~ap_sync_load_value41_U0_ap_ready);
    assign proc_11_output_sync_blk[12] = 1'b0;
    assign proc_dep_vld_vec_11[12] = dl_detect_out ? proc_dep_vld_vec_11_reg[12] : (proc_11_data_FIFO_blk[12] | proc_11_data_PIPO_blk[12] | proc_11_start_FIFO_blk[12] | proc_11_TLF_FIFO_blk[12] | proc_11_input_sync_blk[12] | proc_11_output_sync_blk[12]);
    assign proc_11_data_FIFO_blk[13] = 1'b0;
    assign proc_11_data_PIPO_blk[13] = 1'b0;
    assign proc_11_start_FIFO_blk[13] = 1'b0;
    assign proc_11_TLF_FIFO_blk[13] = 1'b0;
    assign proc_11_input_sync_blk[13] = 1'b0 | (ap_sync_load_value40_U0_ap_ready & load_value40_U0.ap_idle & ~ap_sync_load_value42_U0_ap_ready);
    assign proc_11_output_sync_blk[13] = 1'b0;
    assign proc_dep_vld_vec_11[13] = dl_detect_out ? proc_dep_vld_vec_11_reg[13] : (proc_11_data_FIFO_blk[13] | proc_11_data_PIPO_blk[13] | proc_11_start_FIFO_blk[13] | proc_11_TLF_FIFO_blk[13] | proc_11_input_sync_blk[13] | proc_11_output_sync_blk[13]);
    assign proc_11_data_FIFO_blk[14] = 1'b0;
    assign proc_11_data_PIPO_blk[14] = 1'b0;
    assign proc_11_start_FIFO_blk[14] = 1'b0;
    assign proc_11_TLF_FIFO_blk[14] = 1'b0;
    assign proc_11_input_sync_blk[14] = 1'b0 | (ap_sync_load_value40_U0_ap_ready & load_value40_U0.ap_idle & ~ap_sync_load_value43_U0_ap_ready);
    assign proc_11_output_sync_blk[14] = 1'b0;
    assign proc_dep_vld_vec_11[14] = dl_detect_out ? proc_dep_vld_vec_11_reg[14] : (proc_11_data_FIFO_blk[14] | proc_11_data_PIPO_blk[14] | proc_11_start_FIFO_blk[14] | proc_11_TLF_FIFO_blk[14] | proc_11_input_sync_blk[14] | proc_11_output_sync_blk[14]);
    assign proc_11_data_FIFO_blk[15] = 1'b0;
    assign proc_11_data_PIPO_blk[15] = 1'b0;
    assign proc_11_start_FIFO_blk[15] = 1'b0;
    assign proc_11_TLF_FIFO_blk[15] = 1'b0;
    assign proc_11_input_sync_blk[15] = 1'b0 | (ap_sync_load_value40_U0_ap_ready & load_value40_U0.ap_idle & ~ap_sync_load_value44_U0_ap_ready);
    assign proc_11_output_sync_blk[15] = 1'b0;
    assign proc_dep_vld_vec_11[15] = dl_detect_out ? proc_dep_vld_vec_11_reg[15] : (proc_11_data_FIFO_blk[15] | proc_11_data_PIPO_blk[15] | proc_11_start_FIFO_blk[15] | proc_11_TLF_FIFO_blk[15] | proc_11_input_sync_blk[15] | proc_11_output_sync_blk[15]);
    assign proc_11_data_FIFO_blk[16] = 1'b0;
    assign proc_11_data_PIPO_blk[16] = 1'b0;
    assign proc_11_start_FIFO_blk[16] = 1'b0;
    assign proc_11_TLF_FIFO_blk[16] = 1'b0;
    assign proc_11_input_sync_blk[16] = 1'b0 | (ap_sync_load_value40_U0_ap_ready & load_value40_U0.ap_idle & ~ap_sync_load_value45_U0_ap_ready);
    assign proc_11_output_sync_blk[16] = 1'b0;
    assign proc_dep_vld_vec_11[16] = dl_detect_out ? proc_dep_vld_vec_11_reg[16] : (proc_11_data_FIFO_blk[16] | proc_11_data_PIPO_blk[16] | proc_11_start_FIFO_blk[16] | proc_11_TLF_FIFO_blk[16] | proc_11_input_sync_blk[16] | proc_11_output_sync_blk[16]);
    assign proc_11_data_FIFO_blk[17] = 1'b0;
    assign proc_11_data_PIPO_blk[17] = 1'b0;
    assign proc_11_start_FIFO_blk[17] = 1'b0;
    assign proc_11_TLF_FIFO_blk[17] = 1'b0;
    assign proc_11_input_sync_blk[17] = 1'b0 | (ap_sync_load_value40_U0_ap_ready & load_value40_U0.ap_idle & ~ap_sync_load_value46_U0_ap_ready);
    assign proc_11_output_sync_blk[17] = 1'b0;
    assign proc_dep_vld_vec_11[17] = dl_detect_out ? proc_dep_vld_vec_11_reg[17] : (proc_11_data_FIFO_blk[17] | proc_11_data_PIPO_blk[17] | proc_11_start_FIFO_blk[17] | proc_11_TLF_FIFO_blk[17] | proc_11_input_sync_blk[17] | proc_11_output_sync_blk[17]);
    assign proc_11_data_FIFO_blk[18] = 1'b0;
    assign proc_11_data_PIPO_blk[18] = 1'b0;
    assign proc_11_start_FIFO_blk[18] = 1'b0;
    assign proc_11_TLF_FIFO_blk[18] = 1'b0;
    assign proc_11_input_sync_blk[18] = 1'b0 | (ap_sync_load_value40_U0_ap_ready & load_value40_U0.ap_idle & ~ap_sync_load_value47_U0_ap_ready);
    assign proc_11_output_sync_blk[18] = 1'b0;
    assign proc_dep_vld_vec_11[18] = dl_detect_out ? proc_dep_vld_vec_11_reg[18] : (proc_11_data_FIFO_blk[18] | proc_11_data_PIPO_blk[18] | proc_11_start_FIFO_blk[18] | proc_11_TLF_FIFO_blk[18] | proc_11_input_sync_blk[18] | proc_11_output_sync_blk[18]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_11_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_11_reg <= proc_dep_vld_vec_11;
        end
    end
    assign in_chan_dep_vld_vec_11[0] = dep_chan_vld_0_11;
    assign in_chan_dep_data_vec_11[34 : 0] = dep_chan_data_0_11;
    assign token_in_vec_11[0] = token_0_11;
    assign in_chan_dep_vld_vec_11[1] = dep_chan_vld_1_11;
    assign in_chan_dep_data_vec_11[69 : 35] = dep_chan_data_1_11;
    assign token_in_vec_11[1] = token_1_11;
    assign in_chan_dep_vld_vec_11[2] = dep_chan_vld_2_11;
    assign in_chan_dep_data_vec_11[104 : 70] = dep_chan_data_2_11;
    assign token_in_vec_11[2] = token_2_11;
    assign in_chan_dep_vld_vec_11[3] = dep_chan_vld_3_11;
    assign in_chan_dep_data_vec_11[139 : 105] = dep_chan_data_3_11;
    assign token_in_vec_11[3] = token_3_11;
    assign in_chan_dep_vld_vec_11[4] = dep_chan_vld_4_11;
    assign in_chan_dep_data_vec_11[174 : 140] = dep_chan_data_4_11;
    assign token_in_vec_11[4] = token_4_11;
    assign in_chan_dep_vld_vec_11[5] = dep_chan_vld_5_11;
    assign in_chan_dep_data_vec_11[209 : 175] = dep_chan_data_5_11;
    assign token_in_vec_11[5] = token_5_11;
    assign in_chan_dep_vld_vec_11[6] = dep_chan_vld_6_11;
    assign in_chan_dep_data_vec_11[244 : 210] = dep_chan_data_6_11;
    assign token_in_vec_11[6] = token_6_11;
    assign in_chan_dep_vld_vec_11[7] = dep_chan_vld_7_11;
    assign in_chan_dep_data_vec_11[279 : 245] = dep_chan_data_7_11;
    assign token_in_vec_11[7] = token_7_11;
    assign in_chan_dep_vld_vec_11[8] = dep_chan_vld_8_11;
    assign in_chan_dep_data_vec_11[314 : 280] = dep_chan_data_8_11;
    assign token_in_vec_11[8] = token_8_11;
    assign in_chan_dep_vld_vec_11[9] = dep_chan_vld_9_11;
    assign in_chan_dep_data_vec_11[349 : 315] = dep_chan_data_9_11;
    assign token_in_vec_11[9] = token_9_11;
    assign in_chan_dep_vld_vec_11[10] = dep_chan_vld_10_11;
    assign in_chan_dep_data_vec_11[384 : 350] = dep_chan_data_10_11;
    assign token_in_vec_11[10] = token_10_11;
    assign in_chan_dep_vld_vec_11[11] = dep_chan_vld_12_11;
    assign in_chan_dep_data_vec_11[419 : 385] = dep_chan_data_12_11;
    assign token_in_vec_11[11] = token_12_11;
    assign in_chan_dep_vld_vec_11[12] = dep_chan_vld_13_11;
    assign in_chan_dep_data_vec_11[454 : 420] = dep_chan_data_13_11;
    assign token_in_vec_11[12] = token_13_11;
    assign in_chan_dep_vld_vec_11[13] = dep_chan_vld_14_11;
    assign in_chan_dep_data_vec_11[489 : 455] = dep_chan_data_14_11;
    assign token_in_vec_11[13] = token_14_11;
    assign in_chan_dep_vld_vec_11[14] = dep_chan_vld_15_11;
    assign in_chan_dep_data_vec_11[524 : 490] = dep_chan_data_15_11;
    assign token_in_vec_11[14] = token_15_11;
    assign in_chan_dep_vld_vec_11[15] = dep_chan_vld_16_11;
    assign in_chan_dep_data_vec_11[559 : 525] = dep_chan_data_16_11;
    assign token_in_vec_11[15] = token_16_11;
    assign in_chan_dep_vld_vec_11[16] = dep_chan_vld_17_11;
    assign in_chan_dep_data_vec_11[594 : 560] = dep_chan_data_17_11;
    assign token_in_vec_11[16] = token_17_11;
    assign in_chan_dep_vld_vec_11[17] = dep_chan_vld_18_11;
    assign in_chan_dep_data_vec_11[629 : 595] = dep_chan_data_18_11;
    assign token_in_vec_11[17] = token_18_11;
    assign in_chan_dep_vld_vec_11[18] = dep_chan_vld_27_11;
    assign in_chan_dep_data_vec_11[664 : 630] = dep_chan_data_27_11;
    assign token_in_vec_11[18] = token_27_11;
    assign dep_chan_vld_11_0 = out_chan_dep_vld_vec_11[0];
    assign dep_chan_data_11_0 = out_chan_dep_data_11;
    assign token_11_0 = token_out_vec_11[0];
    assign dep_chan_vld_11_2 = out_chan_dep_vld_vec_11[1];
    assign dep_chan_data_11_2 = out_chan_dep_data_11;
    assign token_11_2 = token_out_vec_11[1];
    assign dep_chan_vld_11_27 = out_chan_dep_vld_vec_11[2];
    assign dep_chan_data_11_27 = out_chan_dep_data_11;
    assign token_11_27 = token_out_vec_11[2];
    assign dep_chan_vld_11_1 = out_chan_dep_vld_vec_11[3];
    assign dep_chan_data_11_1 = out_chan_dep_data_11;
    assign token_11_1 = token_out_vec_11[3];
    assign dep_chan_vld_11_3 = out_chan_dep_vld_vec_11[4];
    assign dep_chan_data_11_3 = out_chan_dep_data_11;
    assign token_11_3 = token_out_vec_11[4];
    assign dep_chan_vld_11_4 = out_chan_dep_vld_vec_11[5];
    assign dep_chan_data_11_4 = out_chan_dep_data_11;
    assign token_11_4 = token_out_vec_11[5];
    assign dep_chan_vld_11_5 = out_chan_dep_vld_vec_11[6];
    assign dep_chan_data_11_5 = out_chan_dep_data_11;
    assign token_11_5 = token_out_vec_11[6];
    assign dep_chan_vld_11_6 = out_chan_dep_vld_vec_11[7];
    assign dep_chan_data_11_6 = out_chan_dep_data_11;
    assign token_11_6 = token_out_vec_11[7];
    assign dep_chan_vld_11_7 = out_chan_dep_vld_vec_11[8];
    assign dep_chan_data_11_7 = out_chan_dep_data_11;
    assign token_11_7 = token_out_vec_11[8];
    assign dep_chan_vld_11_8 = out_chan_dep_vld_vec_11[9];
    assign dep_chan_data_11_8 = out_chan_dep_data_11;
    assign token_11_8 = token_out_vec_11[9];
    assign dep_chan_vld_11_9 = out_chan_dep_vld_vec_11[10];
    assign dep_chan_data_11_9 = out_chan_dep_data_11;
    assign token_11_9 = token_out_vec_11[10];
    assign dep_chan_vld_11_10 = out_chan_dep_vld_vec_11[11];
    assign dep_chan_data_11_10 = out_chan_dep_data_11;
    assign token_11_10 = token_out_vec_11[11];
    assign dep_chan_vld_11_12 = out_chan_dep_vld_vec_11[12];
    assign dep_chan_data_11_12 = out_chan_dep_data_11;
    assign token_11_12 = token_out_vec_11[12];
    assign dep_chan_vld_11_13 = out_chan_dep_vld_vec_11[13];
    assign dep_chan_data_11_13 = out_chan_dep_data_11;
    assign token_11_13 = token_out_vec_11[13];
    assign dep_chan_vld_11_14 = out_chan_dep_vld_vec_11[14];
    assign dep_chan_data_11_14 = out_chan_dep_data_11;
    assign token_11_14 = token_out_vec_11[14];
    assign dep_chan_vld_11_15 = out_chan_dep_vld_vec_11[15];
    assign dep_chan_data_11_15 = out_chan_dep_data_11;
    assign token_11_15 = token_out_vec_11[15];
    assign dep_chan_vld_11_16 = out_chan_dep_vld_vec_11[16];
    assign dep_chan_data_11_16 = out_chan_dep_data_11;
    assign token_11_16 = token_out_vec_11[16];
    assign dep_chan_vld_11_17 = out_chan_dep_vld_vec_11[17];
    assign dep_chan_data_11_17 = out_chan_dep_data_11;
    assign token_11_17 = token_out_vec_11[17];
    assign dep_chan_vld_11_18 = out_chan_dep_vld_vec_11[18];
    assign dep_chan_data_11_18 = out_chan_dep_data_11;
    assign token_11_18 = token_out_vec_11[18];

    // Process: load_value41_U0
    kernel_pr_hls_deadlock_detect_unit #(35, 12, 19, 19) kernel_pr_hls_deadlock_detect_unit_12 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_12),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_12),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_12),
        .token_in_vec(token_in_vec_12),
        .dl_detect_in(dl_detect_out),
        .origin(origin[12]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_12),
        .out_chan_dep_data(out_chan_dep_data_12),
        .token_out_vec(token_out_vec_12),
        .dl_detect_out(dl_in_vec[12]));

    assign proc_12_data_FIFO_blk[0] = 1'b0 | (~load_value41_U0.value_r_blk_n);
    assign proc_12_data_PIPO_blk[0] = 1'b0;
    assign proc_12_start_FIFO_blk[0] = 1'b0;
    assign proc_12_TLF_FIFO_blk[0] = 1'b0;
    assign proc_12_input_sync_blk[0] = 1'b0 | (ap_sync_load_value41_U0_ap_ready & load_value41_U0.ap_idle & ~ap_sync_kernel_pr_entry98_U0_ap_ready);
    assign proc_12_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_12[0] = dl_detect_out ? proc_dep_vld_vec_12_reg[0] : (proc_12_data_FIFO_blk[0] | proc_12_data_PIPO_blk[0] | proc_12_start_FIFO_blk[0] | proc_12_TLF_FIFO_blk[0] | proc_12_input_sync_blk[0] | proc_12_output_sync_blk[0]);
    assign proc_12_data_FIFO_blk[1] = 1'b0 | (~load_value41_U0.bipedge_size_blk_n) | (~load_value41_U0.bipedge_stream_V_V9_blk_n);
    assign proc_12_data_PIPO_blk[1] = 1'b0;
    assign proc_12_start_FIFO_blk[1] = 1'b0;
    assign proc_12_TLF_FIFO_blk[1] = 1'b0;
    assign proc_12_input_sync_blk[1] = 1'b0 | (ap_sync_load_value41_U0_ap_ready & load_value41_U0.ap_idle & ~ap_sync_load_bipedge31_U0_ap_ready);
    assign proc_12_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_12[1] = dl_detect_out ? proc_dep_vld_vec_12_reg[1] : (proc_12_data_FIFO_blk[1] | proc_12_data_PIPO_blk[1] | proc_12_start_FIFO_blk[1] | proc_12_TLF_FIFO_blk[1] | proc_12_input_sync_blk[1] | proc_12_output_sync_blk[1]);
    assign proc_12_data_FIFO_blk[2] = 1'b0 | (~load_value41_U0.value_stream_V_V24_blk_n);
    assign proc_12_data_PIPO_blk[2] = 1'b0;
    assign proc_12_start_FIFO_blk[2] = 1'b0;
    assign proc_12_TLF_FIFO_blk[2] = 1'b0;
    assign proc_12_input_sync_blk[2] = 1'b0;
    assign proc_12_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_12[2] = dl_detect_out ? proc_dep_vld_vec_12_reg[2] : (proc_12_data_FIFO_blk[2] | proc_12_data_PIPO_blk[2] | proc_12_start_FIFO_blk[2] | proc_12_TLF_FIFO_blk[2] | proc_12_input_sync_blk[2] | proc_12_output_sync_blk[2]);
    assign proc_12_data_FIFO_blk[3] = 1'b0;
    assign proc_12_data_PIPO_blk[3] = 1'b0;
    assign proc_12_start_FIFO_blk[3] = 1'b0;
    assign proc_12_TLF_FIFO_blk[3] = 1'b0;
    assign proc_12_input_sync_blk[3] = 1'b0 | (ap_sync_load_value41_U0_ap_ready & load_value41_U0.ap_idle & ~ap_sync_load_bipedge30_U0_ap_ready);
    assign proc_12_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_12[3] = dl_detect_out ? proc_dep_vld_vec_12_reg[3] : (proc_12_data_FIFO_blk[3] | proc_12_data_PIPO_blk[3] | proc_12_start_FIFO_blk[3] | proc_12_TLF_FIFO_blk[3] | proc_12_input_sync_blk[3] | proc_12_output_sync_blk[3]);
    assign proc_12_data_FIFO_blk[4] = 1'b0;
    assign proc_12_data_PIPO_blk[4] = 1'b0;
    assign proc_12_start_FIFO_blk[4] = 1'b0;
    assign proc_12_TLF_FIFO_blk[4] = 1'b0;
    assign proc_12_input_sync_blk[4] = 1'b0 | (ap_sync_load_value41_U0_ap_ready & load_value41_U0.ap_idle & ~ap_sync_load_value32_U0_ap_ready);
    assign proc_12_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_12[4] = dl_detect_out ? proc_dep_vld_vec_12_reg[4] : (proc_12_data_FIFO_blk[4] | proc_12_data_PIPO_blk[4] | proc_12_start_FIFO_blk[4] | proc_12_TLF_FIFO_blk[4] | proc_12_input_sync_blk[4] | proc_12_output_sync_blk[4]);
    assign proc_12_data_FIFO_blk[5] = 1'b0;
    assign proc_12_data_PIPO_blk[5] = 1'b0;
    assign proc_12_start_FIFO_blk[5] = 1'b0;
    assign proc_12_TLF_FIFO_blk[5] = 1'b0;
    assign proc_12_input_sync_blk[5] = 1'b0 | (ap_sync_load_value41_U0_ap_ready & load_value41_U0.ap_idle & ~ap_sync_load_value33_U0_ap_ready);
    assign proc_12_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_12[5] = dl_detect_out ? proc_dep_vld_vec_12_reg[5] : (proc_12_data_FIFO_blk[5] | proc_12_data_PIPO_blk[5] | proc_12_start_FIFO_blk[5] | proc_12_TLF_FIFO_blk[5] | proc_12_input_sync_blk[5] | proc_12_output_sync_blk[5]);
    assign proc_12_data_FIFO_blk[6] = 1'b0;
    assign proc_12_data_PIPO_blk[6] = 1'b0;
    assign proc_12_start_FIFO_blk[6] = 1'b0;
    assign proc_12_TLF_FIFO_blk[6] = 1'b0;
    assign proc_12_input_sync_blk[6] = 1'b0 | (ap_sync_load_value41_U0_ap_ready & load_value41_U0.ap_idle & ~ap_sync_load_value34_U0_ap_ready);
    assign proc_12_output_sync_blk[6] = 1'b0;
    assign proc_dep_vld_vec_12[6] = dl_detect_out ? proc_dep_vld_vec_12_reg[6] : (proc_12_data_FIFO_blk[6] | proc_12_data_PIPO_blk[6] | proc_12_start_FIFO_blk[6] | proc_12_TLF_FIFO_blk[6] | proc_12_input_sync_blk[6] | proc_12_output_sync_blk[6]);
    assign proc_12_data_FIFO_blk[7] = 1'b0;
    assign proc_12_data_PIPO_blk[7] = 1'b0;
    assign proc_12_start_FIFO_blk[7] = 1'b0;
    assign proc_12_TLF_FIFO_blk[7] = 1'b0;
    assign proc_12_input_sync_blk[7] = 1'b0 | (ap_sync_load_value41_U0_ap_ready & load_value41_U0.ap_idle & ~ap_sync_load_value35_U0_ap_ready);
    assign proc_12_output_sync_blk[7] = 1'b0;
    assign proc_dep_vld_vec_12[7] = dl_detect_out ? proc_dep_vld_vec_12_reg[7] : (proc_12_data_FIFO_blk[7] | proc_12_data_PIPO_blk[7] | proc_12_start_FIFO_blk[7] | proc_12_TLF_FIFO_blk[7] | proc_12_input_sync_blk[7] | proc_12_output_sync_blk[7]);
    assign proc_12_data_FIFO_blk[8] = 1'b0;
    assign proc_12_data_PIPO_blk[8] = 1'b0;
    assign proc_12_start_FIFO_blk[8] = 1'b0;
    assign proc_12_TLF_FIFO_blk[8] = 1'b0;
    assign proc_12_input_sync_blk[8] = 1'b0 | (ap_sync_load_value41_U0_ap_ready & load_value41_U0.ap_idle & ~ap_sync_load_value36_U0_ap_ready);
    assign proc_12_output_sync_blk[8] = 1'b0;
    assign proc_dep_vld_vec_12[8] = dl_detect_out ? proc_dep_vld_vec_12_reg[8] : (proc_12_data_FIFO_blk[8] | proc_12_data_PIPO_blk[8] | proc_12_start_FIFO_blk[8] | proc_12_TLF_FIFO_blk[8] | proc_12_input_sync_blk[8] | proc_12_output_sync_blk[8]);
    assign proc_12_data_FIFO_blk[9] = 1'b0;
    assign proc_12_data_PIPO_blk[9] = 1'b0;
    assign proc_12_start_FIFO_blk[9] = 1'b0;
    assign proc_12_TLF_FIFO_blk[9] = 1'b0;
    assign proc_12_input_sync_blk[9] = 1'b0 | (ap_sync_load_value41_U0_ap_ready & load_value41_U0.ap_idle & ~ap_sync_load_value37_U0_ap_ready);
    assign proc_12_output_sync_blk[9] = 1'b0;
    assign proc_dep_vld_vec_12[9] = dl_detect_out ? proc_dep_vld_vec_12_reg[9] : (proc_12_data_FIFO_blk[9] | proc_12_data_PIPO_blk[9] | proc_12_start_FIFO_blk[9] | proc_12_TLF_FIFO_blk[9] | proc_12_input_sync_blk[9] | proc_12_output_sync_blk[9]);
    assign proc_12_data_FIFO_blk[10] = 1'b0;
    assign proc_12_data_PIPO_blk[10] = 1'b0;
    assign proc_12_start_FIFO_blk[10] = 1'b0;
    assign proc_12_TLF_FIFO_blk[10] = 1'b0;
    assign proc_12_input_sync_blk[10] = 1'b0 | (ap_sync_load_value41_U0_ap_ready & load_value41_U0.ap_idle & ~ap_sync_load_value38_U0_ap_ready);
    assign proc_12_output_sync_blk[10] = 1'b0;
    assign proc_dep_vld_vec_12[10] = dl_detect_out ? proc_dep_vld_vec_12_reg[10] : (proc_12_data_FIFO_blk[10] | proc_12_data_PIPO_blk[10] | proc_12_start_FIFO_blk[10] | proc_12_TLF_FIFO_blk[10] | proc_12_input_sync_blk[10] | proc_12_output_sync_blk[10]);
    assign proc_12_data_FIFO_blk[11] = 1'b0;
    assign proc_12_data_PIPO_blk[11] = 1'b0;
    assign proc_12_start_FIFO_blk[11] = 1'b0;
    assign proc_12_TLF_FIFO_blk[11] = 1'b0;
    assign proc_12_input_sync_blk[11] = 1'b0 | (ap_sync_load_value41_U0_ap_ready & load_value41_U0.ap_idle & ~ap_sync_load_value39_U0_ap_ready);
    assign proc_12_output_sync_blk[11] = 1'b0;
    assign proc_dep_vld_vec_12[11] = dl_detect_out ? proc_dep_vld_vec_12_reg[11] : (proc_12_data_FIFO_blk[11] | proc_12_data_PIPO_blk[11] | proc_12_start_FIFO_blk[11] | proc_12_TLF_FIFO_blk[11] | proc_12_input_sync_blk[11] | proc_12_output_sync_blk[11]);
    assign proc_12_data_FIFO_blk[12] = 1'b0;
    assign proc_12_data_PIPO_blk[12] = 1'b0;
    assign proc_12_start_FIFO_blk[12] = 1'b0;
    assign proc_12_TLF_FIFO_blk[12] = 1'b0;
    assign proc_12_input_sync_blk[12] = 1'b0 | (ap_sync_load_value41_U0_ap_ready & load_value41_U0.ap_idle & ~ap_sync_load_value40_U0_ap_ready);
    assign proc_12_output_sync_blk[12] = 1'b0;
    assign proc_dep_vld_vec_12[12] = dl_detect_out ? proc_dep_vld_vec_12_reg[12] : (proc_12_data_FIFO_blk[12] | proc_12_data_PIPO_blk[12] | proc_12_start_FIFO_blk[12] | proc_12_TLF_FIFO_blk[12] | proc_12_input_sync_blk[12] | proc_12_output_sync_blk[12]);
    assign proc_12_data_FIFO_blk[13] = 1'b0;
    assign proc_12_data_PIPO_blk[13] = 1'b0;
    assign proc_12_start_FIFO_blk[13] = 1'b0;
    assign proc_12_TLF_FIFO_blk[13] = 1'b0;
    assign proc_12_input_sync_blk[13] = 1'b0 | (ap_sync_load_value41_U0_ap_ready & load_value41_U0.ap_idle & ~ap_sync_load_value42_U0_ap_ready);
    assign proc_12_output_sync_blk[13] = 1'b0;
    assign proc_dep_vld_vec_12[13] = dl_detect_out ? proc_dep_vld_vec_12_reg[13] : (proc_12_data_FIFO_blk[13] | proc_12_data_PIPO_blk[13] | proc_12_start_FIFO_blk[13] | proc_12_TLF_FIFO_blk[13] | proc_12_input_sync_blk[13] | proc_12_output_sync_blk[13]);
    assign proc_12_data_FIFO_blk[14] = 1'b0;
    assign proc_12_data_PIPO_blk[14] = 1'b0;
    assign proc_12_start_FIFO_blk[14] = 1'b0;
    assign proc_12_TLF_FIFO_blk[14] = 1'b0;
    assign proc_12_input_sync_blk[14] = 1'b0 | (ap_sync_load_value41_U0_ap_ready & load_value41_U0.ap_idle & ~ap_sync_load_value43_U0_ap_ready);
    assign proc_12_output_sync_blk[14] = 1'b0;
    assign proc_dep_vld_vec_12[14] = dl_detect_out ? proc_dep_vld_vec_12_reg[14] : (proc_12_data_FIFO_blk[14] | proc_12_data_PIPO_blk[14] | proc_12_start_FIFO_blk[14] | proc_12_TLF_FIFO_blk[14] | proc_12_input_sync_blk[14] | proc_12_output_sync_blk[14]);
    assign proc_12_data_FIFO_blk[15] = 1'b0;
    assign proc_12_data_PIPO_blk[15] = 1'b0;
    assign proc_12_start_FIFO_blk[15] = 1'b0;
    assign proc_12_TLF_FIFO_blk[15] = 1'b0;
    assign proc_12_input_sync_blk[15] = 1'b0 | (ap_sync_load_value41_U0_ap_ready & load_value41_U0.ap_idle & ~ap_sync_load_value44_U0_ap_ready);
    assign proc_12_output_sync_blk[15] = 1'b0;
    assign proc_dep_vld_vec_12[15] = dl_detect_out ? proc_dep_vld_vec_12_reg[15] : (proc_12_data_FIFO_blk[15] | proc_12_data_PIPO_blk[15] | proc_12_start_FIFO_blk[15] | proc_12_TLF_FIFO_blk[15] | proc_12_input_sync_blk[15] | proc_12_output_sync_blk[15]);
    assign proc_12_data_FIFO_blk[16] = 1'b0;
    assign proc_12_data_PIPO_blk[16] = 1'b0;
    assign proc_12_start_FIFO_blk[16] = 1'b0;
    assign proc_12_TLF_FIFO_blk[16] = 1'b0;
    assign proc_12_input_sync_blk[16] = 1'b0 | (ap_sync_load_value41_U0_ap_ready & load_value41_U0.ap_idle & ~ap_sync_load_value45_U0_ap_ready);
    assign proc_12_output_sync_blk[16] = 1'b0;
    assign proc_dep_vld_vec_12[16] = dl_detect_out ? proc_dep_vld_vec_12_reg[16] : (proc_12_data_FIFO_blk[16] | proc_12_data_PIPO_blk[16] | proc_12_start_FIFO_blk[16] | proc_12_TLF_FIFO_blk[16] | proc_12_input_sync_blk[16] | proc_12_output_sync_blk[16]);
    assign proc_12_data_FIFO_blk[17] = 1'b0;
    assign proc_12_data_PIPO_blk[17] = 1'b0;
    assign proc_12_start_FIFO_blk[17] = 1'b0;
    assign proc_12_TLF_FIFO_blk[17] = 1'b0;
    assign proc_12_input_sync_blk[17] = 1'b0 | (ap_sync_load_value41_U0_ap_ready & load_value41_U0.ap_idle & ~ap_sync_load_value46_U0_ap_ready);
    assign proc_12_output_sync_blk[17] = 1'b0;
    assign proc_dep_vld_vec_12[17] = dl_detect_out ? proc_dep_vld_vec_12_reg[17] : (proc_12_data_FIFO_blk[17] | proc_12_data_PIPO_blk[17] | proc_12_start_FIFO_blk[17] | proc_12_TLF_FIFO_blk[17] | proc_12_input_sync_blk[17] | proc_12_output_sync_blk[17]);
    assign proc_12_data_FIFO_blk[18] = 1'b0;
    assign proc_12_data_PIPO_blk[18] = 1'b0;
    assign proc_12_start_FIFO_blk[18] = 1'b0;
    assign proc_12_TLF_FIFO_blk[18] = 1'b0;
    assign proc_12_input_sync_blk[18] = 1'b0 | (ap_sync_load_value41_U0_ap_ready & load_value41_U0.ap_idle & ~ap_sync_load_value47_U0_ap_ready);
    assign proc_12_output_sync_blk[18] = 1'b0;
    assign proc_dep_vld_vec_12[18] = dl_detect_out ? proc_dep_vld_vec_12_reg[18] : (proc_12_data_FIFO_blk[18] | proc_12_data_PIPO_blk[18] | proc_12_start_FIFO_blk[18] | proc_12_TLF_FIFO_blk[18] | proc_12_input_sync_blk[18] | proc_12_output_sync_blk[18]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_12_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_12_reg <= proc_dep_vld_vec_12;
        end
    end
    assign in_chan_dep_vld_vec_12[0] = dep_chan_vld_0_12;
    assign in_chan_dep_data_vec_12[34 : 0] = dep_chan_data_0_12;
    assign token_in_vec_12[0] = token_0_12;
    assign in_chan_dep_vld_vec_12[1] = dep_chan_vld_1_12;
    assign in_chan_dep_data_vec_12[69 : 35] = dep_chan_data_1_12;
    assign token_in_vec_12[1] = token_1_12;
    assign in_chan_dep_vld_vec_12[2] = dep_chan_vld_2_12;
    assign in_chan_dep_data_vec_12[104 : 70] = dep_chan_data_2_12;
    assign token_in_vec_12[2] = token_2_12;
    assign in_chan_dep_vld_vec_12[3] = dep_chan_vld_3_12;
    assign in_chan_dep_data_vec_12[139 : 105] = dep_chan_data_3_12;
    assign token_in_vec_12[3] = token_3_12;
    assign in_chan_dep_vld_vec_12[4] = dep_chan_vld_4_12;
    assign in_chan_dep_data_vec_12[174 : 140] = dep_chan_data_4_12;
    assign token_in_vec_12[4] = token_4_12;
    assign in_chan_dep_vld_vec_12[5] = dep_chan_vld_5_12;
    assign in_chan_dep_data_vec_12[209 : 175] = dep_chan_data_5_12;
    assign token_in_vec_12[5] = token_5_12;
    assign in_chan_dep_vld_vec_12[6] = dep_chan_vld_6_12;
    assign in_chan_dep_data_vec_12[244 : 210] = dep_chan_data_6_12;
    assign token_in_vec_12[6] = token_6_12;
    assign in_chan_dep_vld_vec_12[7] = dep_chan_vld_7_12;
    assign in_chan_dep_data_vec_12[279 : 245] = dep_chan_data_7_12;
    assign token_in_vec_12[7] = token_7_12;
    assign in_chan_dep_vld_vec_12[8] = dep_chan_vld_8_12;
    assign in_chan_dep_data_vec_12[314 : 280] = dep_chan_data_8_12;
    assign token_in_vec_12[8] = token_8_12;
    assign in_chan_dep_vld_vec_12[9] = dep_chan_vld_9_12;
    assign in_chan_dep_data_vec_12[349 : 315] = dep_chan_data_9_12;
    assign token_in_vec_12[9] = token_9_12;
    assign in_chan_dep_vld_vec_12[10] = dep_chan_vld_10_12;
    assign in_chan_dep_data_vec_12[384 : 350] = dep_chan_data_10_12;
    assign token_in_vec_12[10] = token_10_12;
    assign in_chan_dep_vld_vec_12[11] = dep_chan_vld_11_12;
    assign in_chan_dep_data_vec_12[419 : 385] = dep_chan_data_11_12;
    assign token_in_vec_12[11] = token_11_12;
    assign in_chan_dep_vld_vec_12[12] = dep_chan_vld_13_12;
    assign in_chan_dep_data_vec_12[454 : 420] = dep_chan_data_13_12;
    assign token_in_vec_12[12] = token_13_12;
    assign in_chan_dep_vld_vec_12[13] = dep_chan_vld_14_12;
    assign in_chan_dep_data_vec_12[489 : 455] = dep_chan_data_14_12;
    assign token_in_vec_12[13] = token_14_12;
    assign in_chan_dep_vld_vec_12[14] = dep_chan_vld_15_12;
    assign in_chan_dep_data_vec_12[524 : 490] = dep_chan_data_15_12;
    assign token_in_vec_12[14] = token_15_12;
    assign in_chan_dep_vld_vec_12[15] = dep_chan_vld_16_12;
    assign in_chan_dep_data_vec_12[559 : 525] = dep_chan_data_16_12;
    assign token_in_vec_12[15] = token_16_12;
    assign in_chan_dep_vld_vec_12[16] = dep_chan_vld_17_12;
    assign in_chan_dep_data_vec_12[594 : 560] = dep_chan_data_17_12;
    assign token_in_vec_12[16] = token_17_12;
    assign in_chan_dep_vld_vec_12[17] = dep_chan_vld_18_12;
    assign in_chan_dep_data_vec_12[629 : 595] = dep_chan_data_18_12;
    assign token_in_vec_12[17] = token_18_12;
    assign in_chan_dep_vld_vec_12[18] = dep_chan_vld_28_12;
    assign in_chan_dep_data_vec_12[664 : 630] = dep_chan_data_28_12;
    assign token_in_vec_12[18] = token_28_12;
    assign dep_chan_vld_12_0 = out_chan_dep_vld_vec_12[0];
    assign dep_chan_data_12_0 = out_chan_dep_data_12;
    assign token_12_0 = token_out_vec_12[0];
    assign dep_chan_vld_12_2 = out_chan_dep_vld_vec_12[1];
    assign dep_chan_data_12_2 = out_chan_dep_data_12;
    assign token_12_2 = token_out_vec_12[1];
    assign dep_chan_vld_12_28 = out_chan_dep_vld_vec_12[2];
    assign dep_chan_data_12_28 = out_chan_dep_data_12;
    assign token_12_28 = token_out_vec_12[2];
    assign dep_chan_vld_12_1 = out_chan_dep_vld_vec_12[3];
    assign dep_chan_data_12_1 = out_chan_dep_data_12;
    assign token_12_1 = token_out_vec_12[3];
    assign dep_chan_vld_12_3 = out_chan_dep_vld_vec_12[4];
    assign dep_chan_data_12_3 = out_chan_dep_data_12;
    assign token_12_3 = token_out_vec_12[4];
    assign dep_chan_vld_12_4 = out_chan_dep_vld_vec_12[5];
    assign dep_chan_data_12_4 = out_chan_dep_data_12;
    assign token_12_4 = token_out_vec_12[5];
    assign dep_chan_vld_12_5 = out_chan_dep_vld_vec_12[6];
    assign dep_chan_data_12_5 = out_chan_dep_data_12;
    assign token_12_5 = token_out_vec_12[6];
    assign dep_chan_vld_12_6 = out_chan_dep_vld_vec_12[7];
    assign dep_chan_data_12_6 = out_chan_dep_data_12;
    assign token_12_6 = token_out_vec_12[7];
    assign dep_chan_vld_12_7 = out_chan_dep_vld_vec_12[8];
    assign dep_chan_data_12_7 = out_chan_dep_data_12;
    assign token_12_7 = token_out_vec_12[8];
    assign dep_chan_vld_12_8 = out_chan_dep_vld_vec_12[9];
    assign dep_chan_data_12_8 = out_chan_dep_data_12;
    assign token_12_8 = token_out_vec_12[9];
    assign dep_chan_vld_12_9 = out_chan_dep_vld_vec_12[10];
    assign dep_chan_data_12_9 = out_chan_dep_data_12;
    assign token_12_9 = token_out_vec_12[10];
    assign dep_chan_vld_12_10 = out_chan_dep_vld_vec_12[11];
    assign dep_chan_data_12_10 = out_chan_dep_data_12;
    assign token_12_10 = token_out_vec_12[11];
    assign dep_chan_vld_12_11 = out_chan_dep_vld_vec_12[12];
    assign dep_chan_data_12_11 = out_chan_dep_data_12;
    assign token_12_11 = token_out_vec_12[12];
    assign dep_chan_vld_12_13 = out_chan_dep_vld_vec_12[13];
    assign dep_chan_data_12_13 = out_chan_dep_data_12;
    assign token_12_13 = token_out_vec_12[13];
    assign dep_chan_vld_12_14 = out_chan_dep_vld_vec_12[14];
    assign dep_chan_data_12_14 = out_chan_dep_data_12;
    assign token_12_14 = token_out_vec_12[14];
    assign dep_chan_vld_12_15 = out_chan_dep_vld_vec_12[15];
    assign dep_chan_data_12_15 = out_chan_dep_data_12;
    assign token_12_15 = token_out_vec_12[15];
    assign dep_chan_vld_12_16 = out_chan_dep_vld_vec_12[16];
    assign dep_chan_data_12_16 = out_chan_dep_data_12;
    assign token_12_16 = token_out_vec_12[16];
    assign dep_chan_vld_12_17 = out_chan_dep_vld_vec_12[17];
    assign dep_chan_data_12_17 = out_chan_dep_data_12;
    assign token_12_17 = token_out_vec_12[17];
    assign dep_chan_vld_12_18 = out_chan_dep_vld_vec_12[18];
    assign dep_chan_data_12_18 = out_chan_dep_data_12;
    assign token_12_18 = token_out_vec_12[18];

    // Process: load_value42_U0
    kernel_pr_hls_deadlock_detect_unit #(35, 13, 19, 19) kernel_pr_hls_deadlock_detect_unit_13 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_13),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_13),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_13),
        .token_in_vec(token_in_vec_13),
        .dl_detect_in(dl_detect_out),
        .origin(origin[13]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_13),
        .out_chan_dep_data(out_chan_dep_data_13),
        .token_out_vec(token_out_vec_13),
        .dl_detect_out(dl_in_vec[13]));

    assign proc_13_data_FIFO_blk[0] = 1'b0 | (~load_value42_U0.value_r_blk_n);
    assign proc_13_data_PIPO_blk[0] = 1'b0;
    assign proc_13_start_FIFO_blk[0] = 1'b0;
    assign proc_13_TLF_FIFO_blk[0] = 1'b0;
    assign proc_13_input_sync_blk[0] = 1'b0 | (ap_sync_load_value42_U0_ap_ready & load_value42_U0.ap_idle & ~ap_sync_kernel_pr_entry98_U0_ap_ready);
    assign proc_13_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_13[0] = dl_detect_out ? proc_dep_vld_vec_13_reg[0] : (proc_13_data_FIFO_blk[0] | proc_13_data_PIPO_blk[0] | proc_13_start_FIFO_blk[0] | proc_13_TLF_FIFO_blk[0] | proc_13_input_sync_blk[0] | proc_13_output_sync_blk[0]);
    assign proc_13_data_FIFO_blk[1] = 1'b0 | (~load_value42_U0.bipedge_size_blk_n) | (~load_value42_U0.bipedge_stream_V_V10_blk_n);
    assign proc_13_data_PIPO_blk[1] = 1'b0;
    assign proc_13_start_FIFO_blk[1] = 1'b0;
    assign proc_13_TLF_FIFO_blk[1] = 1'b0;
    assign proc_13_input_sync_blk[1] = 1'b0 | (ap_sync_load_value42_U0_ap_ready & load_value42_U0.ap_idle & ~ap_sync_load_bipedge31_U0_ap_ready);
    assign proc_13_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_13[1] = dl_detect_out ? proc_dep_vld_vec_13_reg[1] : (proc_13_data_FIFO_blk[1] | proc_13_data_PIPO_blk[1] | proc_13_start_FIFO_blk[1] | proc_13_TLF_FIFO_blk[1] | proc_13_input_sync_blk[1] | proc_13_output_sync_blk[1]);
    assign proc_13_data_FIFO_blk[2] = 1'b0 | (~load_value42_U0.value_stream_V_V25_blk_n);
    assign proc_13_data_PIPO_blk[2] = 1'b0;
    assign proc_13_start_FIFO_blk[2] = 1'b0;
    assign proc_13_TLF_FIFO_blk[2] = 1'b0;
    assign proc_13_input_sync_blk[2] = 1'b0;
    assign proc_13_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_13[2] = dl_detect_out ? proc_dep_vld_vec_13_reg[2] : (proc_13_data_FIFO_blk[2] | proc_13_data_PIPO_blk[2] | proc_13_start_FIFO_blk[2] | proc_13_TLF_FIFO_blk[2] | proc_13_input_sync_blk[2] | proc_13_output_sync_blk[2]);
    assign proc_13_data_FIFO_blk[3] = 1'b0;
    assign proc_13_data_PIPO_blk[3] = 1'b0;
    assign proc_13_start_FIFO_blk[3] = 1'b0;
    assign proc_13_TLF_FIFO_blk[3] = 1'b0;
    assign proc_13_input_sync_blk[3] = 1'b0 | (ap_sync_load_value42_U0_ap_ready & load_value42_U0.ap_idle & ~ap_sync_load_bipedge30_U0_ap_ready);
    assign proc_13_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_13[3] = dl_detect_out ? proc_dep_vld_vec_13_reg[3] : (proc_13_data_FIFO_blk[3] | proc_13_data_PIPO_blk[3] | proc_13_start_FIFO_blk[3] | proc_13_TLF_FIFO_blk[3] | proc_13_input_sync_blk[3] | proc_13_output_sync_blk[3]);
    assign proc_13_data_FIFO_blk[4] = 1'b0;
    assign proc_13_data_PIPO_blk[4] = 1'b0;
    assign proc_13_start_FIFO_blk[4] = 1'b0;
    assign proc_13_TLF_FIFO_blk[4] = 1'b0;
    assign proc_13_input_sync_blk[4] = 1'b0 | (ap_sync_load_value42_U0_ap_ready & load_value42_U0.ap_idle & ~ap_sync_load_value32_U0_ap_ready);
    assign proc_13_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_13[4] = dl_detect_out ? proc_dep_vld_vec_13_reg[4] : (proc_13_data_FIFO_blk[4] | proc_13_data_PIPO_blk[4] | proc_13_start_FIFO_blk[4] | proc_13_TLF_FIFO_blk[4] | proc_13_input_sync_blk[4] | proc_13_output_sync_blk[4]);
    assign proc_13_data_FIFO_blk[5] = 1'b0;
    assign proc_13_data_PIPO_blk[5] = 1'b0;
    assign proc_13_start_FIFO_blk[5] = 1'b0;
    assign proc_13_TLF_FIFO_blk[5] = 1'b0;
    assign proc_13_input_sync_blk[5] = 1'b0 | (ap_sync_load_value42_U0_ap_ready & load_value42_U0.ap_idle & ~ap_sync_load_value33_U0_ap_ready);
    assign proc_13_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_13[5] = dl_detect_out ? proc_dep_vld_vec_13_reg[5] : (proc_13_data_FIFO_blk[5] | proc_13_data_PIPO_blk[5] | proc_13_start_FIFO_blk[5] | proc_13_TLF_FIFO_blk[5] | proc_13_input_sync_blk[5] | proc_13_output_sync_blk[5]);
    assign proc_13_data_FIFO_blk[6] = 1'b0;
    assign proc_13_data_PIPO_blk[6] = 1'b0;
    assign proc_13_start_FIFO_blk[6] = 1'b0;
    assign proc_13_TLF_FIFO_blk[6] = 1'b0;
    assign proc_13_input_sync_blk[6] = 1'b0 | (ap_sync_load_value42_U0_ap_ready & load_value42_U0.ap_idle & ~ap_sync_load_value34_U0_ap_ready);
    assign proc_13_output_sync_blk[6] = 1'b0;
    assign proc_dep_vld_vec_13[6] = dl_detect_out ? proc_dep_vld_vec_13_reg[6] : (proc_13_data_FIFO_blk[6] | proc_13_data_PIPO_blk[6] | proc_13_start_FIFO_blk[6] | proc_13_TLF_FIFO_blk[6] | proc_13_input_sync_blk[6] | proc_13_output_sync_blk[6]);
    assign proc_13_data_FIFO_blk[7] = 1'b0;
    assign proc_13_data_PIPO_blk[7] = 1'b0;
    assign proc_13_start_FIFO_blk[7] = 1'b0;
    assign proc_13_TLF_FIFO_blk[7] = 1'b0;
    assign proc_13_input_sync_blk[7] = 1'b0 | (ap_sync_load_value42_U0_ap_ready & load_value42_U0.ap_idle & ~ap_sync_load_value35_U0_ap_ready);
    assign proc_13_output_sync_blk[7] = 1'b0;
    assign proc_dep_vld_vec_13[7] = dl_detect_out ? proc_dep_vld_vec_13_reg[7] : (proc_13_data_FIFO_blk[7] | proc_13_data_PIPO_blk[7] | proc_13_start_FIFO_blk[7] | proc_13_TLF_FIFO_blk[7] | proc_13_input_sync_blk[7] | proc_13_output_sync_blk[7]);
    assign proc_13_data_FIFO_blk[8] = 1'b0;
    assign proc_13_data_PIPO_blk[8] = 1'b0;
    assign proc_13_start_FIFO_blk[8] = 1'b0;
    assign proc_13_TLF_FIFO_blk[8] = 1'b0;
    assign proc_13_input_sync_blk[8] = 1'b0 | (ap_sync_load_value42_U0_ap_ready & load_value42_U0.ap_idle & ~ap_sync_load_value36_U0_ap_ready);
    assign proc_13_output_sync_blk[8] = 1'b0;
    assign proc_dep_vld_vec_13[8] = dl_detect_out ? proc_dep_vld_vec_13_reg[8] : (proc_13_data_FIFO_blk[8] | proc_13_data_PIPO_blk[8] | proc_13_start_FIFO_blk[8] | proc_13_TLF_FIFO_blk[8] | proc_13_input_sync_blk[8] | proc_13_output_sync_blk[8]);
    assign proc_13_data_FIFO_blk[9] = 1'b0;
    assign proc_13_data_PIPO_blk[9] = 1'b0;
    assign proc_13_start_FIFO_blk[9] = 1'b0;
    assign proc_13_TLF_FIFO_blk[9] = 1'b0;
    assign proc_13_input_sync_blk[9] = 1'b0 | (ap_sync_load_value42_U0_ap_ready & load_value42_U0.ap_idle & ~ap_sync_load_value37_U0_ap_ready);
    assign proc_13_output_sync_blk[9] = 1'b0;
    assign proc_dep_vld_vec_13[9] = dl_detect_out ? proc_dep_vld_vec_13_reg[9] : (proc_13_data_FIFO_blk[9] | proc_13_data_PIPO_blk[9] | proc_13_start_FIFO_blk[9] | proc_13_TLF_FIFO_blk[9] | proc_13_input_sync_blk[9] | proc_13_output_sync_blk[9]);
    assign proc_13_data_FIFO_blk[10] = 1'b0;
    assign proc_13_data_PIPO_blk[10] = 1'b0;
    assign proc_13_start_FIFO_blk[10] = 1'b0;
    assign proc_13_TLF_FIFO_blk[10] = 1'b0;
    assign proc_13_input_sync_blk[10] = 1'b0 | (ap_sync_load_value42_U0_ap_ready & load_value42_U0.ap_idle & ~ap_sync_load_value38_U0_ap_ready);
    assign proc_13_output_sync_blk[10] = 1'b0;
    assign proc_dep_vld_vec_13[10] = dl_detect_out ? proc_dep_vld_vec_13_reg[10] : (proc_13_data_FIFO_blk[10] | proc_13_data_PIPO_blk[10] | proc_13_start_FIFO_blk[10] | proc_13_TLF_FIFO_blk[10] | proc_13_input_sync_blk[10] | proc_13_output_sync_blk[10]);
    assign proc_13_data_FIFO_blk[11] = 1'b0;
    assign proc_13_data_PIPO_blk[11] = 1'b0;
    assign proc_13_start_FIFO_blk[11] = 1'b0;
    assign proc_13_TLF_FIFO_blk[11] = 1'b0;
    assign proc_13_input_sync_blk[11] = 1'b0 | (ap_sync_load_value42_U0_ap_ready & load_value42_U0.ap_idle & ~ap_sync_load_value39_U0_ap_ready);
    assign proc_13_output_sync_blk[11] = 1'b0;
    assign proc_dep_vld_vec_13[11] = dl_detect_out ? proc_dep_vld_vec_13_reg[11] : (proc_13_data_FIFO_blk[11] | proc_13_data_PIPO_blk[11] | proc_13_start_FIFO_blk[11] | proc_13_TLF_FIFO_blk[11] | proc_13_input_sync_blk[11] | proc_13_output_sync_blk[11]);
    assign proc_13_data_FIFO_blk[12] = 1'b0;
    assign proc_13_data_PIPO_blk[12] = 1'b0;
    assign proc_13_start_FIFO_blk[12] = 1'b0;
    assign proc_13_TLF_FIFO_blk[12] = 1'b0;
    assign proc_13_input_sync_blk[12] = 1'b0 | (ap_sync_load_value42_U0_ap_ready & load_value42_U0.ap_idle & ~ap_sync_load_value40_U0_ap_ready);
    assign proc_13_output_sync_blk[12] = 1'b0;
    assign proc_dep_vld_vec_13[12] = dl_detect_out ? proc_dep_vld_vec_13_reg[12] : (proc_13_data_FIFO_blk[12] | proc_13_data_PIPO_blk[12] | proc_13_start_FIFO_blk[12] | proc_13_TLF_FIFO_blk[12] | proc_13_input_sync_blk[12] | proc_13_output_sync_blk[12]);
    assign proc_13_data_FIFO_blk[13] = 1'b0;
    assign proc_13_data_PIPO_blk[13] = 1'b0;
    assign proc_13_start_FIFO_blk[13] = 1'b0;
    assign proc_13_TLF_FIFO_blk[13] = 1'b0;
    assign proc_13_input_sync_blk[13] = 1'b0 | (ap_sync_load_value42_U0_ap_ready & load_value42_U0.ap_idle & ~ap_sync_load_value41_U0_ap_ready);
    assign proc_13_output_sync_blk[13] = 1'b0;
    assign proc_dep_vld_vec_13[13] = dl_detect_out ? proc_dep_vld_vec_13_reg[13] : (proc_13_data_FIFO_blk[13] | proc_13_data_PIPO_blk[13] | proc_13_start_FIFO_blk[13] | proc_13_TLF_FIFO_blk[13] | proc_13_input_sync_blk[13] | proc_13_output_sync_blk[13]);
    assign proc_13_data_FIFO_blk[14] = 1'b0;
    assign proc_13_data_PIPO_blk[14] = 1'b0;
    assign proc_13_start_FIFO_blk[14] = 1'b0;
    assign proc_13_TLF_FIFO_blk[14] = 1'b0;
    assign proc_13_input_sync_blk[14] = 1'b0 | (ap_sync_load_value42_U0_ap_ready & load_value42_U0.ap_idle & ~ap_sync_load_value43_U0_ap_ready);
    assign proc_13_output_sync_blk[14] = 1'b0;
    assign proc_dep_vld_vec_13[14] = dl_detect_out ? proc_dep_vld_vec_13_reg[14] : (proc_13_data_FIFO_blk[14] | proc_13_data_PIPO_blk[14] | proc_13_start_FIFO_blk[14] | proc_13_TLF_FIFO_blk[14] | proc_13_input_sync_blk[14] | proc_13_output_sync_blk[14]);
    assign proc_13_data_FIFO_blk[15] = 1'b0;
    assign proc_13_data_PIPO_blk[15] = 1'b0;
    assign proc_13_start_FIFO_blk[15] = 1'b0;
    assign proc_13_TLF_FIFO_blk[15] = 1'b0;
    assign proc_13_input_sync_blk[15] = 1'b0 | (ap_sync_load_value42_U0_ap_ready & load_value42_U0.ap_idle & ~ap_sync_load_value44_U0_ap_ready);
    assign proc_13_output_sync_blk[15] = 1'b0;
    assign proc_dep_vld_vec_13[15] = dl_detect_out ? proc_dep_vld_vec_13_reg[15] : (proc_13_data_FIFO_blk[15] | proc_13_data_PIPO_blk[15] | proc_13_start_FIFO_blk[15] | proc_13_TLF_FIFO_blk[15] | proc_13_input_sync_blk[15] | proc_13_output_sync_blk[15]);
    assign proc_13_data_FIFO_blk[16] = 1'b0;
    assign proc_13_data_PIPO_blk[16] = 1'b0;
    assign proc_13_start_FIFO_blk[16] = 1'b0;
    assign proc_13_TLF_FIFO_blk[16] = 1'b0;
    assign proc_13_input_sync_blk[16] = 1'b0 | (ap_sync_load_value42_U0_ap_ready & load_value42_U0.ap_idle & ~ap_sync_load_value45_U0_ap_ready);
    assign proc_13_output_sync_blk[16] = 1'b0;
    assign proc_dep_vld_vec_13[16] = dl_detect_out ? proc_dep_vld_vec_13_reg[16] : (proc_13_data_FIFO_blk[16] | proc_13_data_PIPO_blk[16] | proc_13_start_FIFO_blk[16] | proc_13_TLF_FIFO_blk[16] | proc_13_input_sync_blk[16] | proc_13_output_sync_blk[16]);
    assign proc_13_data_FIFO_blk[17] = 1'b0;
    assign proc_13_data_PIPO_blk[17] = 1'b0;
    assign proc_13_start_FIFO_blk[17] = 1'b0;
    assign proc_13_TLF_FIFO_blk[17] = 1'b0;
    assign proc_13_input_sync_blk[17] = 1'b0 | (ap_sync_load_value42_U0_ap_ready & load_value42_U0.ap_idle & ~ap_sync_load_value46_U0_ap_ready);
    assign proc_13_output_sync_blk[17] = 1'b0;
    assign proc_dep_vld_vec_13[17] = dl_detect_out ? proc_dep_vld_vec_13_reg[17] : (proc_13_data_FIFO_blk[17] | proc_13_data_PIPO_blk[17] | proc_13_start_FIFO_blk[17] | proc_13_TLF_FIFO_blk[17] | proc_13_input_sync_blk[17] | proc_13_output_sync_blk[17]);
    assign proc_13_data_FIFO_blk[18] = 1'b0;
    assign proc_13_data_PIPO_blk[18] = 1'b0;
    assign proc_13_start_FIFO_blk[18] = 1'b0;
    assign proc_13_TLF_FIFO_blk[18] = 1'b0;
    assign proc_13_input_sync_blk[18] = 1'b0 | (ap_sync_load_value42_U0_ap_ready & load_value42_U0.ap_idle & ~ap_sync_load_value47_U0_ap_ready);
    assign proc_13_output_sync_blk[18] = 1'b0;
    assign proc_dep_vld_vec_13[18] = dl_detect_out ? proc_dep_vld_vec_13_reg[18] : (proc_13_data_FIFO_blk[18] | proc_13_data_PIPO_blk[18] | proc_13_start_FIFO_blk[18] | proc_13_TLF_FIFO_blk[18] | proc_13_input_sync_blk[18] | proc_13_output_sync_blk[18]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_13_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_13_reg <= proc_dep_vld_vec_13;
        end
    end
    assign in_chan_dep_vld_vec_13[0] = dep_chan_vld_0_13;
    assign in_chan_dep_data_vec_13[34 : 0] = dep_chan_data_0_13;
    assign token_in_vec_13[0] = token_0_13;
    assign in_chan_dep_vld_vec_13[1] = dep_chan_vld_1_13;
    assign in_chan_dep_data_vec_13[69 : 35] = dep_chan_data_1_13;
    assign token_in_vec_13[1] = token_1_13;
    assign in_chan_dep_vld_vec_13[2] = dep_chan_vld_2_13;
    assign in_chan_dep_data_vec_13[104 : 70] = dep_chan_data_2_13;
    assign token_in_vec_13[2] = token_2_13;
    assign in_chan_dep_vld_vec_13[3] = dep_chan_vld_3_13;
    assign in_chan_dep_data_vec_13[139 : 105] = dep_chan_data_3_13;
    assign token_in_vec_13[3] = token_3_13;
    assign in_chan_dep_vld_vec_13[4] = dep_chan_vld_4_13;
    assign in_chan_dep_data_vec_13[174 : 140] = dep_chan_data_4_13;
    assign token_in_vec_13[4] = token_4_13;
    assign in_chan_dep_vld_vec_13[5] = dep_chan_vld_5_13;
    assign in_chan_dep_data_vec_13[209 : 175] = dep_chan_data_5_13;
    assign token_in_vec_13[5] = token_5_13;
    assign in_chan_dep_vld_vec_13[6] = dep_chan_vld_6_13;
    assign in_chan_dep_data_vec_13[244 : 210] = dep_chan_data_6_13;
    assign token_in_vec_13[6] = token_6_13;
    assign in_chan_dep_vld_vec_13[7] = dep_chan_vld_7_13;
    assign in_chan_dep_data_vec_13[279 : 245] = dep_chan_data_7_13;
    assign token_in_vec_13[7] = token_7_13;
    assign in_chan_dep_vld_vec_13[8] = dep_chan_vld_8_13;
    assign in_chan_dep_data_vec_13[314 : 280] = dep_chan_data_8_13;
    assign token_in_vec_13[8] = token_8_13;
    assign in_chan_dep_vld_vec_13[9] = dep_chan_vld_9_13;
    assign in_chan_dep_data_vec_13[349 : 315] = dep_chan_data_9_13;
    assign token_in_vec_13[9] = token_9_13;
    assign in_chan_dep_vld_vec_13[10] = dep_chan_vld_10_13;
    assign in_chan_dep_data_vec_13[384 : 350] = dep_chan_data_10_13;
    assign token_in_vec_13[10] = token_10_13;
    assign in_chan_dep_vld_vec_13[11] = dep_chan_vld_11_13;
    assign in_chan_dep_data_vec_13[419 : 385] = dep_chan_data_11_13;
    assign token_in_vec_13[11] = token_11_13;
    assign in_chan_dep_vld_vec_13[12] = dep_chan_vld_12_13;
    assign in_chan_dep_data_vec_13[454 : 420] = dep_chan_data_12_13;
    assign token_in_vec_13[12] = token_12_13;
    assign in_chan_dep_vld_vec_13[13] = dep_chan_vld_14_13;
    assign in_chan_dep_data_vec_13[489 : 455] = dep_chan_data_14_13;
    assign token_in_vec_13[13] = token_14_13;
    assign in_chan_dep_vld_vec_13[14] = dep_chan_vld_15_13;
    assign in_chan_dep_data_vec_13[524 : 490] = dep_chan_data_15_13;
    assign token_in_vec_13[14] = token_15_13;
    assign in_chan_dep_vld_vec_13[15] = dep_chan_vld_16_13;
    assign in_chan_dep_data_vec_13[559 : 525] = dep_chan_data_16_13;
    assign token_in_vec_13[15] = token_16_13;
    assign in_chan_dep_vld_vec_13[16] = dep_chan_vld_17_13;
    assign in_chan_dep_data_vec_13[594 : 560] = dep_chan_data_17_13;
    assign token_in_vec_13[16] = token_17_13;
    assign in_chan_dep_vld_vec_13[17] = dep_chan_vld_18_13;
    assign in_chan_dep_data_vec_13[629 : 595] = dep_chan_data_18_13;
    assign token_in_vec_13[17] = token_18_13;
    assign in_chan_dep_vld_vec_13[18] = dep_chan_vld_29_13;
    assign in_chan_dep_data_vec_13[664 : 630] = dep_chan_data_29_13;
    assign token_in_vec_13[18] = token_29_13;
    assign dep_chan_vld_13_0 = out_chan_dep_vld_vec_13[0];
    assign dep_chan_data_13_0 = out_chan_dep_data_13;
    assign token_13_0 = token_out_vec_13[0];
    assign dep_chan_vld_13_2 = out_chan_dep_vld_vec_13[1];
    assign dep_chan_data_13_2 = out_chan_dep_data_13;
    assign token_13_2 = token_out_vec_13[1];
    assign dep_chan_vld_13_29 = out_chan_dep_vld_vec_13[2];
    assign dep_chan_data_13_29 = out_chan_dep_data_13;
    assign token_13_29 = token_out_vec_13[2];
    assign dep_chan_vld_13_1 = out_chan_dep_vld_vec_13[3];
    assign dep_chan_data_13_1 = out_chan_dep_data_13;
    assign token_13_1 = token_out_vec_13[3];
    assign dep_chan_vld_13_3 = out_chan_dep_vld_vec_13[4];
    assign dep_chan_data_13_3 = out_chan_dep_data_13;
    assign token_13_3 = token_out_vec_13[4];
    assign dep_chan_vld_13_4 = out_chan_dep_vld_vec_13[5];
    assign dep_chan_data_13_4 = out_chan_dep_data_13;
    assign token_13_4 = token_out_vec_13[5];
    assign dep_chan_vld_13_5 = out_chan_dep_vld_vec_13[6];
    assign dep_chan_data_13_5 = out_chan_dep_data_13;
    assign token_13_5 = token_out_vec_13[6];
    assign dep_chan_vld_13_6 = out_chan_dep_vld_vec_13[7];
    assign dep_chan_data_13_6 = out_chan_dep_data_13;
    assign token_13_6 = token_out_vec_13[7];
    assign dep_chan_vld_13_7 = out_chan_dep_vld_vec_13[8];
    assign dep_chan_data_13_7 = out_chan_dep_data_13;
    assign token_13_7 = token_out_vec_13[8];
    assign dep_chan_vld_13_8 = out_chan_dep_vld_vec_13[9];
    assign dep_chan_data_13_8 = out_chan_dep_data_13;
    assign token_13_8 = token_out_vec_13[9];
    assign dep_chan_vld_13_9 = out_chan_dep_vld_vec_13[10];
    assign dep_chan_data_13_9 = out_chan_dep_data_13;
    assign token_13_9 = token_out_vec_13[10];
    assign dep_chan_vld_13_10 = out_chan_dep_vld_vec_13[11];
    assign dep_chan_data_13_10 = out_chan_dep_data_13;
    assign token_13_10 = token_out_vec_13[11];
    assign dep_chan_vld_13_11 = out_chan_dep_vld_vec_13[12];
    assign dep_chan_data_13_11 = out_chan_dep_data_13;
    assign token_13_11 = token_out_vec_13[12];
    assign dep_chan_vld_13_12 = out_chan_dep_vld_vec_13[13];
    assign dep_chan_data_13_12 = out_chan_dep_data_13;
    assign token_13_12 = token_out_vec_13[13];
    assign dep_chan_vld_13_14 = out_chan_dep_vld_vec_13[14];
    assign dep_chan_data_13_14 = out_chan_dep_data_13;
    assign token_13_14 = token_out_vec_13[14];
    assign dep_chan_vld_13_15 = out_chan_dep_vld_vec_13[15];
    assign dep_chan_data_13_15 = out_chan_dep_data_13;
    assign token_13_15 = token_out_vec_13[15];
    assign dep_chan_vld_13_16 = out_chan_dep_vld_vec_13[16];
    assign dep_chan_data_13_16 = out_chan_dep_data_13;
    assign token_13_16 = token_out_vec_13[16];
    assign dep_chan_vld_13_17 = out_chan_dep_vld_vec_13[17];
    assign dep_chan_data_13_17 = out_chan_dep_data_13;
    assign token_13_17 = token_out_vec_13[17];
    assign dep_chan_vld_13_18 = out_chan_dep_vld_vec_13[18];
    assign dep_chan_data_13_18 = out_chan_dep_data_13;
    assign token_13_18 = token_out_vec_13[18];

    // Process: load_value43_U0
    kernel_pr_hls_deadlock_detect_unit #(35, 14, 19, 19) kernel_pr_hls_deadlock_detect_unit_14 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_14),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_14),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_14),
        .token_in_vec(token_in_vec_14),
        .dl_detect_in(dl_detect_out),
        .origin(origin[14]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_14),
        .out_chan_dep_data(out_chan_dep_data_14),
        .token_out_vec(token_out_vec_14),
        .dl_detect_out(dl_in_vec[14]));

    assign proc_14_data_FIFO_blk[0] = 1'b0 | (~load_value43_U0.value_r_blk_n);
    assign proc_14_data_PIPO_blk[0] = 1'b0;
    assign proc_14_start_FIFO_blk[0] = 1'b0;
    assign proc_14_TLF_FIFO_blk[0] = 1'b0;
    assign proc_14_input_sync_blk[0] = 1'b0 | (ap_sync_load_value43_U0_ap_ready & load_value43_U0.ap_idle & ~ap_sync_kernel_pr_entry98_U0_ap_ready);
    assign proc_14_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_14[0] = dl_detect_out ? proc_dep_vld_vec_14_reg[0] : (proc_14_data_FIFO_blk[0] | proc_14_data_PIPO_blk[0] | proc_14_start_FIFO_blk[0] | proc_14_TLF_FIFO_blk[0] | proc_14_input_sync_blk[0] | proc_14_output_sync_blk[0]);
    assign proc_14_data_FIFO_blk[1] = 1'b0 | (~load_value43_U0.bipedge_size_blk_n) | (~load_value43_U0.bipedge_stream_V_V11_blk_n);
    assign proc_14_data_PIPO_blk[1] = 1'b0;
    assign proc_14_start_FIFO_blk[1] = 1'b0;
    assign proc_14_TLF_FIFO_blk[1] = 1'b0;
    assign proc_14_input_sync_blk[1] = 1'b0 | (ap_sync_load_value43_U0_ap_ready & load_value43_U0.ap_idle & ~ap_sync_load_bipedge31_U0_ap_ready);
    assign proc_14_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_14[1] = dl_detect_out ? proc_dep_vld_vec_14_reg[1] : (proc_14_data_FIFO_blk[1] | proc_14_data_PIPO_blk[1] | proc_14_start_FIFO_blk[1] | proc_14_TLF_FIFO_blk[1] | proc_14_input_sync_blk[1] | proc_14_output_sync_blk[1]);
    assign proc_14_data_FIFO_blk[2] = 1'b0 | (~load_value43_U0.value_stream_V_V26_blk_n);
    assign proc_14_data_PIPO_blk[2] = 1'b0;
    assign proc_14_start_FIFO_blk[2] = 1'b0;
    assign proc_14_TLF_FIFO_blk[2] = 1'b0;
    assign proc_14_input_sync_blk[2] = 1'b0;
    assign proc_14_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_14[2] = dl_detect_out ? proc_dep_vld_vec_14_reg[2] : (proc_14_data_FIFO_blk[2] | proc_14_data_PIPO_blk[2] | proc_14_start_FIFO_blk[2] | proc_14_TLF_FIFO_blk[2] | proc_14_input_sync_blk[2] | proc_14_output_sync_blk[2]);
    assign proc_14_data_FIFO_blk[3] = 1'b0;
    assign proc_14_data_PIPO_blk[3] = 1'b0;
    assign proc_14_start_FIFO_blk[3] = 1'b0;
    assign proc_14_TLF_FIFO_blk[3] = 1'b0;
    assign proc_14_input_sync_blk[3] = 1'b0 | (ap_sync_load_value43_U0_ap_ready & load_value43_U0.ap_idle & ~ap_sync_load_bipedge30_U0_ap_ready);
    assign proc_14_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_14[3] = dl_detect_out ? proc_dep_vld_vec_14_reg[3] : (proc_14_data_FIFO_blk[3] | proc_14_data_PIPO_blk[3] | proc_14_start_FIFO_blk[3] | proc_14_TLF_FIFO_blk[3] | proc_14_input_sync_blk[3] | proc_14_output_sync_blk[3]);
    assign proc_14_data_FIFO_blk[4] = 1'b0;
    assign proc_14_data_PIPO_blk[4] = 1'b0;
    assign proc_14_start_FIFO_blk[4] = 1'b0;
    assign proc_14_TLF_FIFO_blk[4] = 1'b0;
    assign proc_14_input_sync_blk[4] = 1'b0 | (ap_sync_load_value43_U0_ap_ready & load_value43_U0.ap_idle & ~ap_sync_load_value32_U0_ap_ready);
    assign proc_14_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_14[4] = dl_detect_out ? proc_dep_vld_vec_14_reg[4] : (proc_14_data_FIFO_blk[4] | proc_14_data_PIPO_blk[4] | proc_14_start_FIFO_blk[4] | proc_14_TLF_FIFO_blk[4] | proc_14_input_sync_blk[4] | proc_14_output_sync_blk[4]);
    assign proc_14_data_FIFO_blk[5] = 1'b0;
    assign proc_14_data_PIPO_blk[5] = 1'b0;
    assign proc_14_start_FIFO_blk[5] = 1'b0;
    assign proc_14_TLF_FIFO_blk[5] = 1'b0;
    assign proc_14_input_sync_blk[5] = 1'b0 | (ap_sync_load_value43_U0_ap_ready & load_value43_U0.ap_idle & ~ap_sync_load_value33_U0_ap_ready);
    assign proc_14_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_14[5] = dl_detect_out ? proc_dep_vld_vec_14_reg[5] : (proc_14_data_FIFO_blk[5] | proc_14_data_PIPO_blk[5] | proc_14_start_FIFO_blk[5] | proc_14_TLF_FIFO_blk[5] | proc_14_input_sync_blk[5] | proc_14_output_sync_blk[5]);
    assign proc_14_data_FIFO_blk[6] = 1'b0;
    assign proc_14_data_PIPO_blk[6] = 1'b0;
    assign proc_14_start_FIFO_blk[6] = 1'b0;
    assign proc_14_TLF_FIFO_blk[6] = 1'b0;
    assign proc_14_input_sync_blk[6] = 1'b0 | (ap_sync_load_value43_U0_ap_ready & load_value43_U0.ap_idle & ~ap_sync_load_value34_U0_ap_ready);
    assign proc_14_output_sync_blk[6] = 1'b0;
    assign proc_dep_vld_vec_14[6] = dl_detect_out ? proc_dep_vld_vec_14_reg[6] : (proc_14_data_FIFO_blk[6] | proc_14_data_PIPO_blk[6] | proc_14_start_FIFO_blk[6] | proc_14_TLF_FIFO_blk[6] | proc_14_input_sync_blk[6] | proc_14_output_sync_blk[6]);
    assign proc_14_data_FIFO_blk[7] = 1'b0;
    assign proc_14_data_PIPO_blk[7] = 1'b0;
    assign proc_14_start_FIFO_blk[7] = 1'b0;
    assign proc_14_TLF_FIFO_blk[7] = 1'b0;
    assign proc_14_input_sync_blk[7] = 1'b0 | (ap_sync_load_value43_U0_ap_ready & load_value43_U0.ap_idle & ~ap_sync_load_value35_U0_ap_ready);
    assign proc_14_output_sync_blk[7] = 1'b0;
    assign proc_dep_vld_vec_14[7] = dl_detect_out ? proc_dep_vld_vec_14_reg[7] : (proc_14_data_FIFO_blk[7] | proc_14_data_PIPO_blk[7] | proc_14_start_FIFO_blk[7] | proc_14_TLF_FIFO_blk[7] | proc_14_input_sync_blk[7] | proc_14_output_sync_blk[7]);
    assign proc_14_data_FIFO_blk[8] = 1'b0;
    assign proc_14_data_PIPO_blk[8] = 1'b0;
    assign proc_14_start_FIFO_blk[8] = 1'b0;
    assign proc_14_TLF_FIFO_blk[8] = 1'b0;
    assign proc_14_input_sync_blk[8] = 1'b0 | (ap_sync_load_value43_U0_ap_ready & load_value43_U0.ap_idle & ~ap_sync_load_value36_U0_ap_ready);
    assign proc_14_output_sync_blk[8] = 1'b0;
    assign proc_dep_vld_vec_14[8] = dl_detect_out ? proc_dep_vld_vec_14_reg[8] : (proc_14_data_FIFO_blk[8] | proc_14_data_PIPO_blk[8] | proc_14_start_FIFO_blk[8] | proc_14_TLF_FIFO_blk[8] | proc_14_input_sync_blk[8] | proc_14_output_sync_blk[8]);
    assign proc_14_data_FIFO_blk[9] = 1'b0;
    assign proc_14_data_PIPO_blk[9] = 1'b0;
    assign proc_14_start_FIFO_blk[9] = 1'b0;
    assign proc_14_TLF_FIFO_blk[9] = 1'b0;
    assign proc_14_input_sync_blk[9] = 1'b0 | (ap_sync_load_value43_U0_ap_ready & load_value43_U0.ap_idle & ~ap_sync_load_value37_U0_ap_ready);
    assign proc_14_output_sync_blk[9] = 1'b0;
    assign proc_dep_vld_vec_14[9] = dl_detect_out ? proc_dep_vld_vec_14_reg[9] : (proc_14_data_FIFO_blk[9] | proc_14_data_PIPO_blk[9] | proc_14_start_FIFO_blk[9] | proc_14_TLF_FIFO_blk[9] | proc_14_input_sync_blk[9] | proc_14_output_sync_blk[9]);
    assign proc_14_data_FIFO_blk[10] = 1'b0;
    assign proc_14_data_PIPO_blk[10] = 1'b0;
    assign proc_14_start_FIFO_blk[10] = 1'b0;
    assign proc_14_TLF_FIFO_blk[10] = 1'b0;
    assign proc_14_input_sync_blk[10] = 1'b0 | (ap_sync_load_value43_U0_ap_ready & load_value43_U0.ap_idle & ~ap_sync_load_value38_U0_ap_ready);
    assign proc_14_output_sync_blk[10] = 1'b0;
    assign proc_dep_vld_vec_14[10] = dl_detect_out ? proc_dep_vld_vec_14_reg[10] : (proc_14_data_FIFO_blk[10] | proc_14_data_PIPO_blk[10] | proc_14_start_FIFO_blk[10] | proc_14_TLF_FIFO_blk[10] | proc_14_input_sync_blk[10] | proc_14_output_sync_blk[10]);
    assign proc_14_data_FIFO_blk[11] = 1'b0;
    assign proc_14_data_PIPO_blk[11] = 1'b0;
    assign proc_14_start_FIFO_blk[11] = 1'b0;
    assign proc_14_TLF_FIFO_blk[11] = 1'b0;
    assign proc_14_input_sync_blk[11] = 1'b0 | (ap_sync_load_value43_U0_ap_ready & load_value43_U0.ap_idle & ~ap_sync_load_value39_U0_ap_ready);
    assign proc_14_output_sync_blk[11] = 1'b0;
    assign proc_dep_vld_vec_14[11] = dl_detect_out ? proc_dep_vld_vec_14_reg[11] : (proc_14_data_FIFO_blk[11] | proc_14_data_PIPO_blk[11] | proc_14_start_FIFO_blk[11] | proc_14_TLF_FIFO_blk[11] | proc_14_input_sync_blk[11] | proc_14_output_sync_blk[11]);
    assign proc_14_data_FIFO_blk[12] = 1'b0;
    assign proc_14_data_PIPO_blk[12] = 1'b0;
    assign proc_14_start_FIFO_blk[12] = 1'b0;
    assign proc_14_TLF_FIFO_blk[12] = 1'b0;
    assign proc_14_input_sync_blk[12] = 1'b0 | (ap_sync_load_value43_U0_ap_ready & load_value43_U0.ap_idle & ~ap_sync_load_value40_U0_ap_ready);
    assign proc_14_output_sync_blk[12] = 1'b0;
    assign proc_dep_vld_vec_14[12] = dl_detect_out ? proc_dep_vld_vec_14_reg[12] : (proc_14_data_FIFO_blk[12] | proc_14_data_PIPO_blk[12] | proc_14_start_FIFO_blk[12] | proc_14_TLF_FIFO_blk[12] | proc_14_input_sync_blk[12] | proc_14_output_sync_blk[12]);
    assign proc_14_data_FIFO_blk[13] = 1'b0;
    assign proc_14_data_PIPO_blk[13] = 1'b0;
    assign proc_14_start_FIFO_blk[13] = 1'b0;
    assign proc_14_TLF_FIFO_blk[13] = 1'b0;
    assign proc_14_input_sync_blk[13] = 1'b0 | (ap_sync_load_value43_U0_ap_ready & load_value43_U0.ap_idle & ~ap_sync_load_value41_U0_ap_ready);
    assign proc_14_output_sync_blk[13] = 1'b0;
    assign proc_dep_vld_vec_14[13] = dl_detect_out ? proc_dep_vld_vec_14_reg[13] : (proc_14_data_FIFO_blk[13] | proc_14_data_PIPO_blk[13] | proc_14_start_FIFO_blk[13] | proc_14_TLF_FIFO_blk[13] | proc_14_input_sync_blk[13] | proc_14_output_sync_blk[13]);
    assign proc_14_data_FIFO_blk[14] = 1'b0;
    assign proc_14_data_PIPO_blk[14] = 1'b0;
    assign proc_14_start_FIFO_blk[14] = 1'b0;
    assign proc_14_TLF_FIFO_blk[14] = 1'b0;
    assign proc_14_input_sync_blk[14] = 1'b0 | (ap_sync_load_value43_U0_ap_ready & load_value43_U0.ap_idle & ~ap_sync_load_value42_U0_ap_ready);
    assign proc_14_output_sync_blk[14] = 1'b0;
    assign proc_dep_vld_vec_14[14] = dl_detect_out ? proc_dep_vld_vec_14_reg[14] : (proc_14_data_FIFO_blk[14] | proc_14_data_PIPO_blk[14] | proc_14_start_FIFO_blk[14] | proc_14_TLF_FIFO_blk[14] | proc_14_input_sync_blk[14] | proc_14_output_sync_blk[14]);
    assign proc_14_data_FIFO_blk[15] = 1'b0;
    assign proc_14_data_PIPO_blk[15] = 1'b0;
    assign proc_14_start_FIFO_blk[15] = 1'b0;
    assign proc_14_TLF_FIFO_blk[15] = 1'b0;
    assign proc_14_input_sync_blk[15] = 1'b0 | (ap_sync_load_value43_U0_ap_ready & load_value43_U0.ap_idle & ~ap_sync_load_value44_U0_ap_ready);
    assign proc_14_output_sync_blk[15] = 1'b0;
    assign proc_dep_vld_vec_14[15] = dl_detect_out ? proc_dep_vld_vec_14_reg[15] : (proc_14_data_FIFO_blk[15] | proc_14_data_PIPO_blk[15] | proc_14_start_FIFO_blk[15] | proc_14_TLF_FIFO_blk[15] | proc_14_input_sync_blk[15] | proc_14_output_sync_blk[15]);
    assign proc_14_data_FIFO_blk[16] = 1'b0;
    assign proc_14_data_PIPO_blk[16] = 1'b0;
    assign proc_14_start_FIFO_blk[16] = 1'b0;
    assign proc_14_TLF_FIFO_blk[16] = 1'b0;
    assign proc_14_input_sync_blk[16] = 1'b0 | (ap_sync_load_value43_U0_ap_ready & load_value43_U0.ap_idle & ~ap_sync_load_value45_U0_ap_ready);
    assign proc_14_output_sync_blk[16] = 1'b0;
    assign proc_dep_vld_vec_14[16] = dl_detect_out ? proc_dep_vld_vec_14_reg[16] : (proc_14_data_FIFO_blk[16] | proc_14_data_PIPO_blk[16] | proc_14_start_FIFO_blk[16] | proc_14_TLF_FIFO_blk[16] | proc_14_input_sync_blk[16] | proc_14_output_sync_blk[16]);
    assign proc_14_data_FIFO_blk[17] = 1'b0;
    assign proc_14_data_PIPO_blk[17] = 1'b0;
    assign proc_14_start_FIFO_blk[17] = 1'b0;
    assign proc_14_TLF_FIFO_blk[17] = 1'b0;
    assign proc_14_input_sync_blk[17] = 1'b0 | (ap_sync_load_value43_U0_ap_ready & load_value43_U0.ap_idle & ~ap_sync_load_value46_U0_ap_ready);
    assign proc_14_output_sync_blk[17] = 1'b0;
    assign proc_dep_vld_vec_14[17] = dl_detect_out ? proc_dep_vld_vec_14_reg[17] : (proc_14_data_FIFO_blk[17] | proc_14_data_PIPO_blk[17] | proc_14_start_FIFO_blk[17] | proc_14_TLF_FIFO_blk[17] | proc_14_input_sync_blk[17] | proc_14_output_sync_blk[17]);
    assign proc_14_data_FIFO_blk[18] = 1'b0;
    assign proc_14_data_PIPO_blk[18] = 1'b0;
    assign proc_14_start_FIFO_blk[18] = 1'b0;
    assign proc_14_TLF_FIFO_blk[18] = 1'b0;
    assign proc_14_input_sync_blk[18] = 1'b0 | (ap_sync_load_value43_U0_ap_ready & load_value43_U0.ap_idle & ~ap_sync_load_value47_U0_ap_ready);
    assign proc_14_output_sync_blk[18] = 1'b0;
    assign proc_dep_vld_vec_14[18] = dl_detect_out ? proc_dep_vld_vec_14_reg[18] : (proc_14_data_FIFO_blk[18] | proc_14_data_PIPO_blk[18] | proc_14_start_FIFO_blk[18] | proc_14_TLF_FIFO_blk[18] | proc_14_input_sync_blk[18] | proc_14_output_sync_blk[18]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_14_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_14_reg <= proc_dep_vld_vec_14;
        end
    end
    assign in_chan_dep_vld_vec_14[0] = dep_chan_vld_0_14;
    assign in_chan_dep_data_vec_14[34 : 0] = dep_chan_data_0_14;
    assign token_in_vec_14[0] = token_0_14;
    assign in_chan_dep_vld_vec_14[1] = dep_chan_vld_1_14;
    assign in_chan_dep_data_vec_14[69 : 35] = dep_chan_data_1_14;
    assign token_in_vec_14[1] = token_1_14;
    assign in_chan_dep_vld_vec_14[2] = dep_chan_vld_2_14;
    assign in_chan_dep_data_vec_14[104 : 70] = dep_chan_data_2_14;
    assign token_in_vec_14[2] = token_2_14;
    assign in_chan_dep_vld_vec_14[3] = dep_chan_vld_3_14;
    assign in_chan_dep_data_vec_14[139 : 105] = dep_chan_data_3_14;
    assign token_in_vec_14[3] = token_3_14;
    assign in_chan_dep_vld_vec_14[4] = dep_chan_vld_4_14;
    assign in_chan_dep_data_vec_14[174 : 140] = dep_chan_data_4_14;
    assign token_in_vec_14[4] = token_4_14;
    assign in_chan_dep_vld_vec_14[5] = dep_chan_vld_5_14;
    assign in_chan_dep_data_vec_14[209 : 175] = dep_chan_data_5_14;
    assign token_in_vec_14[5] = token_5_14;
    assign in_chan_dep_vld_vec_14[6] = dep_chan_vld_6_14;
    assign in_chan_dep_data_vec_14[244 : 210] = dep_chan_data_6_14;
    assign token_in_vec_14[6] = token_6_14;
    assign in_chan_dep_vld_vec_14[7] = dep_chan_vld_7_14;
    assign in_chan_dep_data_vec_14[279 : 245] = dep_chan_data_7_14;
    assign token_in_vec_14[7] = token_7_14;
    assign in_chan_dep_vld_vec_14[8] = dep_chan_vld_8_14;
    assign in_chan_dep_data_vec_14[314 : 280] = dep_chan_data_8_14;
    assign token_in_vec_14[8] = token_8_14;
    assign in_chan_dep_vld_vec_14[9] = dep_chan_vld_9_14;
    assign in_chan_dep_data_vec_14[349 : 315] = dep_chan_data_9_14;
    assign token_in_vec_14[9] = token_9_14;
    assign in_chan_dep_vld_vec_14[10] = dep_chan_vld_10_14;
    assign in_chan_dep_data_vec_14[384 : 350] = dep_chan_data_10_14;
    assign token_in_vec_14[10] = token_10_14;
    assign in_chan_dep_vld_vec_14[11] = dep_chan_vld_11_14;
    assign in_chan_dep_data_vec_14[419 : 385] = dep_chan_data_11_14;
    assign token_in_vec_14[11] = token_11_14;
    assign in_chan_dep_vld_vec_14[12] = dep_chan_vld_12_14;
    assign in_chan_dep_data_vec_14[454 : 420] = dep_chan_data_12_14;
    assign token_in_vec_14[12] = token_12_14;
    assign in_chan_dep_vld_vec_14[13] = dep_chan_vld_13_14;
    assign in_chan_dep_data_vec_14[489 : 455] = dep_chan_data_13_14;
    assign token_in_vec_14[13] = token_13_14;
    assign in_chan_dep_vld_vec_14[14] = dep_chan_vld_15_14;
    assign in_chan_dep_data_vec_14[524 : 490] = dep_chan_data_15_14;
    assign token_in_vec_14[14] = token_15_14;
    assign in_chan_dep_vld_vec_14[15] = dep_chan_vld_16_14;
    assign in_chan_dep_data_vec_14[559 : 525] = dep_chan_data_16_14;
    assign token_in_vec_14[15] = token_16_14;
    assign in_chan_dep_vld_vec_14[16] = dep_chan_vld_17_14;
    assign in_chan_dep_data_vec_14[594 : 560] = dep_chan_data_17_14;
    assign token_in_vec_14[16] = token_17_14;
    assign in_chan_dep_vld_vec_14[17] = dep_chan_vld_18_14;
    assign in_chan_dep_data_vec_14[629 : 595] = dep_chan_data_18_14;
    assign token_in_vec_14[17] = token_18_14;
    assign in_chan_dep_vld_vec_14[18] = dep_chan_vld_30_14;
    assign in_chan_dep_data_vec_14[664 : 630] = dep_chan_data_30_14;
    assign token_in_vec_14[18] = token_30_14;
    assign dep_chan_vld_14_0 = out_chan_dep_vld_vec_14[0];
    assign dep_chan_data_14_0 = out_chan_dep_data_14;
    assign token_14_0 = token_out_vec_14[0];
    assign dep_chan_vld_14_2 = out_chan_dep_vld_vec_14[1];
    assign dep_chan_data_14_2 = out_chan_dep_data_14;
    assign token_14_2 = token_out_vec_14[1];
    assign dep_chan_vld_14_30 = out_chan_dep_vld_vec_14[2];
    assign dep_chan_data_14_30 = out_chan_dep_data_14;
    assign token_14_30 = token_out_vec_14[2];
    assign dep_chan_vld_14_1 = out_chan_dep_vld_vec_14[3];
    assign dep_chan_data_14_1 = out_chan_dep_data_14;
    assign token_14_1 = token_out_vec_14[3];
    assign dep_chan_vld_14_3 = out_chan_dep_vld_vec_14[4];
    assign dep_chan_data_14_3 = out_chan_dep_data_14;
    assign token_14_3 = token_out_vec_14[4];
    assign dep_chan_vld_14_4 = out_chan_dep_vld_vec_14[5];
    assign dep_chan_data_14_4 = out_chan_dep_data_14;
    assign token_14_4 = token_out_vec_14[5];
    assign dep_chan_vld_14_5 = out_chan_dep_vld_vec_14[6];
    assign dep_chan_data_14_5 = out_chan_dep_data_14;
    assign token_14_5 = token_out_vec_14[6];
    assign dep_chan_vld_14_6 = out_chan_dep_vld_vec_14[7];
    assign dep_chan_data_14_6 = out_chan_dep_data_14;
    assign token_14_6 = token_out_vec_14[7];
    assign dep_chan_vld_14_7 = out_chan_dep_vld_vec_14[8];
    assign dep_chan_data_14_7 = out_chan_dep_data_14;
    assign token_14_7 = token_out_vec_14[8];
    assign dep_chan_vld_14_8 = out_chan_dep_vld_vec_14[9];
    assign dep_chan_data_14_8 = out_chan_dep_data_14;
    assign token_14_8 = token_out_vec_14[9];
    assign dep_chan_vld_14_9 = out_chan_dep_vld_vec_14[10];
    assign dep_chan_data_14_9 = out_chan_dep_data_14;
    assign token_14_9 = token_out_vec_14[10];
    assign dep_chan_vld_14_10 = out_chan_dep_vld_vec_14[11];
    assign dep_chan_data_14_10 = out_chan_dep_data_14;
    assign token_14_10 = token_out_vec_14[11];
    assign dep_chan_vld_14_11 = out_chan_dep_vld_vec_14[12];
    assign dep_chan_data_14_11 = out_chan_dep_data_14;
    assign token_14_11 = token_out_vec_14[12];
    assign dep_chan_vld_14_12 = out_chan_dep_vld_vec_14[13];
    assign dep_chan_data_14_12 = out_chan_dep_data_14;
    assign token_14_12 = token_out_vec_14[13];
    assign dep_chan_vld_14_13 = out_chan_dep_vld_vec_14[14];
    assign dep_chan_data_14_13 = out_chan_dep_data_14;
    assign token_14_13 = token_out_vec_14[14];
    assign dep_chan_vld_14_15 = out_chan_dep_vld_vec_14[15];
    assign dep_chan_data_14_15 = out_chan_dep_data_14;
    assign token_14_15 = token_out_vec_14[15];
    assign dep_chan_vld_14_16 = out_chan_dep_vld_vec_14[16];
    assign dep_chan_data_14_16 = out_chan_dep_data_14;
    assign token_14_16 = token_out_vec_14[16];
    assign dep_chan_vld_14_17 = out_chan_dep_vld_vec_14[17];
    assign dep_chan_data_14_17 = out_chan_dep_data_14;
    assign token_14_17 = token_out_vec_14[17];
    assign dep_chan_vld_14_18 = out_chan_dep_vld_vec_14[18];
    assign dep_chan_data_14_18 = out_chan_dep_data_14;
    assign token_14_18 = token_out_vec_14[18];

    // Process: load_value44_U0
    kernel_pr_hls_deadlock_detect_unit #(35, 15, 19, 19) kernel_pr_hls_deadlock_detect_unit_15 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_15),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_15),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_15),
        .token_in_vec(token_in_vec_15),
        .dl_detect_in(dl_detect_out),
        .origin(origin[15]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_15),
        .out_chan_dep_data(out_chan_dep_data_15),
        .token_out_vec(token_out_vec_15),
        .dl_detect_out(dl_in_vec[15]));

    assign proc_15_data_FIFO_blk[0] = 1'b0 | (~load_value44_U0.value_r_blk_n);
    assign proc_15_data_PIPO_blk[0] = 1'b0;
    assign proc_15_start_FIFO_blk[0] = 1'b0;
    assign proc_15_TLF_FIFO_blk[0] = 1'b0;
    assign proc_15_input_sync_blk[0] = 1'b0 | (ap_sync_load_value44_U0_ap_ready & load_value44_U0.ap_idle & ~ap_sync_kernel_pr_entry98_U0_ap_ready);
    assign proc_15_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_15[0] = dl_detect_out ? proc_dep_vld_vec_15_reg[0] : (proc_15_data_FIFO_blk[0] | proc_15_data_PIPO_blk[0] | proc_15_start_FIFO_blk[0] | proc_15_TLF_FIFO_blk[0] | proc_15_input_sync_blk[0] | proc_15_output_sync_blk[0]);
    assign proc_15_data_FIFO_blk[1] = 1'b0 | (~load_value44_U0.bipedge_size_blk_n) | (~load_value44_U0.bipedge_stream_V_V12_blk_n);
    assign proc_15_data_PIPO_blk[1] = 1'b0;
    assign proc_15_start_FIFO_blk[1] = 1'b0;
    assign proc_15_TLF_FIFO_blk[1] = 1'b0;
    assign proc_15_input_sync_blk[1] = 1'b0 | (ap_sync_load_value44_U0_ap_ready & load_value44_U0.ap_idle & ~ap_sync_load_bipedge31_U0_ap_ready);
    assign proc_15_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_15[1] = dl_detect_out ? proc_dep_vld_vec_15_reg[1] : (proc_15_data_FIFO_blk[1] | proc_15_data_PIPO_blk[1] | proc_15_start_FIFO_blk[1] | proc_15_TLF_FIFO_blk[1] | proc_15_input_sync_blk[1] | proc_15_output_sync_blk[1]);
    assign proc_15_data_FIFO_blk[2] = 1'b0 | (~load_value44_U0.value_stream_V_V27_blk_n);
    assign proc_15_data_PIPO_blk[2] = 1'b0;
    assign proc_15_start_FIFO_blk[2] = 1'b0;
    assign proc_15_TLF_FIFO_blk[2] = 1'b0;
    assign proc_15_input_sync_blk[2] = 1'b0;
    assign proc_15_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_15[2] = dl_detect_out ? proc_dep_vld_vec_15_reg[2] : (proc_15_data_FIFO_blk[2] | proc_15_data_PIPO_blk[2] | proc_15_start_FIFO_blk[2] | proc_15_TLF_FIFO_blk[2] | proc_15_input_sync_blk[2] | proc_15_output_sync_blk[2]);
    assign proc_15_data_FIFO_blk[3] = 1'b0;
    assign proc_15_data_PIPO_blk[3] = 1'b0;
    assign proc_15_start_FIFO_blk[3] = 1'b0;
    assign proc_15_TLF_FIFO_blk[3] = 1'b0;
    assign proc_15_input_sync_blk[3] = 1'b0 | (ap_sync_load_value44_U0_ap_ready & load_value44_U0.ap_idle & ~ap_sync_load_bipedge30_U0_ap_ready);
    assign proc_15_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_15[3] = dl_detect_out ? proc_dep_vld_vec_15_reg[3] : (proc_15_data_FIFO_blk[3] | proc_15_data_PIPO_blk[3] | proc_15_start_FIFO_blk[3] | proc_15_TLF_FIFO_blk[3] | proc_15_input_sync_blk[3] | proc_15_output_sync_blk[3]);
    assign proc_15_data_FIFO_blk[4] = 1'b0;
    assign proc_15_data_PIPO_blk[4] = 1'b0;
    assign proc_15_start_FIFO_blk[4] = 1'b0;
    assign proc_15_TLF_FIFO_blk[4] = 1'b0;
    assign proc_15_input_sync_blk[4] = 1'b0 | (ap_sync_load_value44_U0_ap_ready & load_value44_U0.ap_idle & ~ap_sync_load_value32_U0_ap_ready);
    assign proc_15_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_15[4] = dl_detect_out ? proc_dep_vld_vec_15_reg[4] : (proc_15_data_FIFO_blk[4] | proc_15_data_PIPO_blk[4] | proc_15_start_FIFO_blk[4] | proc_15_TLF_FIFO_blk[4] | proc_15_input_sync_blk[4] | proc_15_output_sync_blk[4]);
    assign proc_15_data_FIFO_blk[5] = 1'b0;
    assign proc_15_data_PIPO_blk[5] = 1'b0;
    assign proc_15_start_FIFO_blk[5] = 1'b0;
    assign proc_15_TLF_FIFO_blk[5] = 1'b0;
    assign proc_15_input_sync_blk[5] = 1'b0 | (ap_sync_load_value44_U0_ap_ready & load_value44_U0.ap_idle & ~ap_sync_load_value33_U0_ap_ready);
    assign proc_15_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_15[5] = dl_detect_out ? proc_dep_vld_vec_15_reg[5] : (proc_15_data_FIFO_blk[5] | proc_15_data_PIPO_blk[5] | proc_15_start_FIFO_blk[5] | proc_15_TLF_FIFO_blk[5] | proc_15_input_sync_blk[5] | proc_15_output_sync_blk[5]);
    assign proc_15_data_FIFO_blk[6] = 1'b0;
    assign proc_15_data_PIPO_blk[6] = 1'b0;
    assign proc_15_start_FIFO_blk[6] = 1'b0;
    assign proc_15_TLF_FIFO_blk[6] = 1'b0;
    assign proc_15_input_sync_blk[6] = 1'b0 | (ap_sync_load_value44_U0_ap_ready & load_value44_U0.ap_idle & ~ap_sync_load_value34_U0_ap_ready);
    assign proc_15_output_sync_blk[6] = 1'b0;
    assign proc_dep_vld_vec_15[6] = dl_detect_out ? proc_dep_vld_vec_15_reg[6] : (proc_15_data_FIFO_blk[6] | proc_15_data_PIPO_blk[6] | proc_15_start_FIFO_blk[6] | proc_15_TLF_FIFO_blk[6] | proc_15_input_sync_blk[6] | proc_15_output_sync_blk[6]);
    assign proc_15_data_FIFO_blk[7] = 1'b0;
    assign proc_15_data_PIPO_blk[7] = 1'b0;
    assign proc_15_start_FIFO_blk[7] = 1'b0;
    assign proc_15_TLF_FIFO_blk[7] = 1'b0;
    assign proc_15_input_sync_blk[7] = 1'b0 | (ap_sync_load_value44_U0_ap_ready & load_value44_U0.ap_idle & ~ap_sync_load_value35_U0_ap_ready);
    assign proc_15_output_sync_blk[7] = 1'b0;
    assign proc_dep_vld_vec_15[7] = dl_detect_out ? proc_dep_vld_vec_15_reg[7] : (proc_15_data_FIFO_blk[7] | proc_15_data_PIPO_blk[7] | proc_15_start_FIFO_blk[7] | proc_15_TLF_FIFO_blk[7] | proc_15_input_sync_blk[7] | proc_15_output_sync_blk[7]);
    assign proc_15_data_FIFO_blk[8] = 1'b0;
    assign proc_15_data_PIPO_blk[8] = 1'b0;
    assign proc_15_start_FIFO_blk[8] = 1'b0;
    assign proc_15_TLF_FIFO_blk[8] = 1'b0;
    assign proc_15_input_sync_blk[8] = 1'b0 | (ap_sync_load_value44_U0_ap_ready & load_value44_U0.ap_idle & ~ap_sync_load_value36_U0_ap_ready);
    assign proc_15_output_sync_blk[8] = 1'b0;
    assign proc_dep_vld_vec_15[8] = dl_detect_out ? proc_dep_vld_vec_15_reg[8] : (proc_15_data_FIFO_blk[8] | proc_15_data_PIPO_blk[8] | proc_15_start_FIFO_blk[8] | proc_15_TLF_FIFO_blk[8] | proc_15_input_sync_blk[8] | proc_15_output_sync_blk[8]);
    assign proc_15_data_FIFO_blk[9] = 1'b0;
    assign proc_15_data_PIPO_blk[9] = 1'b0;
    assign proc_15_start_FIFO_blk[9] = 1'b0;
    assign proc_15_TLF_FIFO_blk[9] = 1'b0;
    assign proc_15_input_sync_blk[9] = 1'b0 | (ap_sync_load_value44_U0_ap_ready & load_value44_U0.ap_idle & ~ap_sync_load_value37_U0_ap_ready);
    assign proc_15_output_sync_blk[9] = 1'b0;
    assign proc_dep_vld_vec_15[9] = dl_detect_out ? proc_dep_vld_vec_15_reg[9] : (proc_15_data_FIFO_blk[9] | proc_15_data_PIPO_blk[9] | proc_15_start_FIFO_blk[9] | proc_15_TLF_FIFO_blk[9] | proc_15_input_sync_blk[9] | proc_15_output_sync_blk[9]);
    assign proc_15_data_FIFO_blk[10] = 1'b0;
    assign proc_15_data_PIPO_blk[10] = 1'b0;
    assign proc_15_start_FIFO_blk[10] = 1'b0;
    assign proc_15_TLF_FIFO_blk[10] = 1'b0;
    assign proc_15_input_sync_blk[10] = 1'b0 | (ap_sync_load_value44_U0_ap_ready & load_value44_U0.ap_idle & ~ap_sync_load_value38_U0_ap_ready);
    assign proc_15_output_sync_blk[10] = 1'b0;
    assign proc_dep_vld_vec_15[10] = dl_detect_out ? proc_dep_vld_vec_15_reg[10] : (proc_15_data_FIFO_blk[10] | proc_15_data_PIPO_blk[10] | proc_15_start_FIFO_blk[10] | proc_15_TLF_FIFO_blk[10] | proc_15_input_sync_blk[10] | proc_15_output_sync_blk[10]);
    assign proc_15_data_FIFO_blk[11] = 1'b0;
    assign proc_15_data_PIPO_blk[11] = 1'b0;
    assign proc_15_start_FIFO_blk[11] = 1'b0;
    assign proc_15_TLF_FIFO_blk[11] = 1'b0;
    assign proc_15_input_sync_blk[11] = 1'b0 | (ap_sync_load_value44_U0_ap_ready & load_value44_U0.ap_idle & ~ap_sync_load_value39_U0_ap_ready);
    assign proc_15_output_sync_blk[11] = 1'b0;
    assign proc_dep_vld_vec_15[11] = dl_detect_out ? proc_dep_vld_vec_15_reg[11] : (proc_15_data_FIFO_blk[11] | proc_15_data_PIPO_blk[11] | proc_15_start_FIFO_blk[11] | proc_15_TLF_FIFO_blk[11] | proc_15_input_sync_blk[11] | proc_15_output_sync_blk[11]);
    assign proc_15_data_FIFO_blk[12] = 1'b0;
    assign proc_15_data_PIPO_blk[12] = 1'b0;
    assign proc_15_start_FIFO_blk[12] = 1'b0;
    assign proc_15_TLF_FIFO_blk[12] = 1'b0;
    assign proc_15_input_sync_blk[12] = 1'b0 | (ap_sync_load_value44_U0_ap_ready & load_value44_U0.ap_idle & ~ap_sync_load_value40_U0_ap_ready);
    assign proc_15_output_sync_blk[12] = 1'b0;
    assign proc_dep_vld_vec_15[12] = dl_detect_out ? proc_dep_vld_vec_15_reg[12] : (proc_15_data_FIFO_blk[12] | proc_15_data_PIPO_blk[12] | proc_15_start_FIFO_blk[12] | proc_15_TLF_FIFO_blk[12] | proc_15_input_sync_blk[12] | proc_15_output_sync_blk[12]);
    assign proc_15_data_FIFO_blk[13] = 1'b0;
    assign proc_15_data_PIPO_blk[13] = 1'b0;
    assign proc_15_start_FIFO_blk[13] = 1'b0;
    assign proc_15_TLF_FIFO_blk[13] = 1'b0;
    assign proc_15_input_sync_blk[13] = 1'b0 | (ap_sync_load_value44_U0_ap_ready & load_value44_U0.ap_idle & ~ap_sync_load_value41_U0_ap_ready);
    assign proc_15_output_sync_blk[13] = 1'b0;
    assign proc_dep_vld_vec_15[13] = dl_detect_out ? proc_dep_vld_vec_15_reg[13] : (proc_15_data_FIFO_blk[13] | proc_15_data_PIPO_blk[13] | proc_15_start_FIFO_blk[13] | proc_15_TLF_FIFO_blk[13] | proc_15_input_sync_blk[13] | proc_15_output_sync_blk[13]);
    assign proc_15_data_FIFO_blk[14] = 1'b0;
    assign proc_15_data_PIPO_blk[14] = 1'b0;
    assign proc_15_start_FIFO_blk[14] = 1'b0;
    assign proc_15_TLF_FIFO_blk[14] = 1'b0;
    assign proc_15_input_sync_blk[14] = 1'b0 | (ap_sync_load_value44_U0_ap_ready & load_value44_U0.ap_idle & ~ap_sync_load_value42_U0_ap_ready);
    assign proc_15_output_sync_blk[14] = 1'b0;
    assign proc_dep_vld_vec_15[14] = dl_detect_out ? proc_dep_vld_vec_15_reg[14] : (proc_15_data_FIFO_blk[14] | proc_15_data_PIPO_blk[14] | proc_15_start_FIFO_blk[14] | proc_15_TLF_FIFO_blk[14] | proc_15_input_sync_blk[14] | proc_15_output_sync_blk[14]);
    assign proc_15_data_FIFO_blk[15] = 1'b0;
    assign proc_15_data_PIPO_blk[15] = 1'b0;
    assign proc_15_start_FIFO_blk[15] = 1'b0;
    assign proc_15_TLF_FIFO_blk[15] = 1'b0;
    assign proc_15_input_sync_blk[15] = 1'b0 | (ap_sync_load_value44_U0_ap_ready & load_value44_U0.ap_idle & ~ap_sync_load_value43_U0_ap_ready);
    assign proc_15_output_sync_blk[15] = 1'b0;
    assign proc_dep_vld_vec_15[15] = dl_detect_out ? proc_dep_vld_vec_15_reg[15] : (proc_15_data_FIFO_blk[15] | proc_15_data_PIPO_blk[15] | proc_15_start_FIFO_blk[15] | proc_15_TLF_FIFO_blk[15] | proc_15_input_sync_blk[15] | proc_15_output_sync_blk[15]);
    assign proc_15_data_FIFO_blk[16] = 1'b0;
    assign proc_15_data_PIPO_blk[16] = 1'b0;
    assign proc_15_start_FIFO_blk[16] = 1'b0;
    assign proc_15_TLF_FIFO_blk[16] = 1'b0;
    assign proc_15_input_sync_blk[16] = 1'b0 | (ap_sync_load_value44_U0_ap_ready & load_value44_U0.ap_idle & ~ap_sync_load_value45_U0_ap_ready);
    assign proc_15_output_sync_blk[16] = 1'b0;
    assign proc_dep_vld_vec_15[16] = dl_detect_out ? proc_dep_vld_vec_15_reg[16] : (proc_15_data_FIFO_blk[16] | proc_15_data_PIPO_blk[16] | proc_15_start_FIFO_blk[16] | proc_15_TLF_FIFO_blk[16] | proc_15_input_sync_blk[16] | proc_15_output_sync_blk[16]);
    assign proc_15_data_FIFO_blk[17] = 1'b0;
    assign proc_15_data_PIPO_blk[17] = 1'b0;
    assign proc_15_start_FIFO_blk[17] = 1'b0;
    assign proc_15_TLF_FIFO_blk[17] = 1'b0;
    assign proc_15_input_sync_blk[17] = 1'b0 | (ap_sync_load_value44_U0_ap_ready & load_value44_U0.ap_idle & ~ap_sync_load_value46_U0_ap_ready);
    assign proc_15_output_sync_blk[17] = 1'b0;
    assign proc_dep_vld_vec_15[17] = dl_detect_out ? proc_dep_vld_vec_15_reg[17] : (proc_15_data_FIFO_blk[17] | proc_15_data_PIPO_blk[17] | proc_15_start_FIFO_blk[17] | proc_15_TLF_FIFO_blk[17] | proc_15_input_sync_blk[17] | proc_15_output_sync_blk[17]);
    assign proc_15_data_FIFO_blk[18] = 1'b0;
    assign proc_15_data_PIPO_blk[18] = 1'b0;
    assign proc_15_start_FIFO_blk[18] = 1'b0;
    assign proc_15_TLF_FIFO_blk[18] = 1'b0;
    assign proc_15_input_sync_blk[18] = 1'b0 | (ap_sync_load_value44_U0_ap_ready & load_value44_U0.ap_idle & ~ap_sync_load_value47_U0_ap_ready);
    assign proc_15_output_sync_blk[18] = 1'b0;
    assign proc_dep_vld_vec_15[18] = dl_detect_out ? proc_dep_vld_vec_15_reg[18] : (proc_15_data_FIFO_blk[18] | proc_15_data_PIPO_blk[18] | proc_15_start_FIFO_blk[18] | proc_15_TLF_FIFO_blk[18] | proc_15_input_sync_blk[18] | proc_15_output_sync_blk[18]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_15_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_15_reg <= proc_dep_vld_vec_15;
        end
    end
    assign in_chan_dep_vld_vec_15[0] = dep_chan_vld_0_15;
    assign in_chan_dep_data_vec_15[34 : 0] = dep_chan_data_0_15;
    assign token_in_vec_15[0] = token_0_15;
    assign in_chan_dep_vld_vec_15[1] = dep_chan_vld_1_15;
    assign in_chan_dep_data_vec_15[69 : 35] = dep_chan_data_1_15;
    assign token_in_vec_15[1] = token_1_15;
    assign in_chan_dep_vld_vec_15[2] = dep_chan_vld_2_15;
    assign in_chan_dep_data_vec_15[104 : 70] = dep_chan_data_2_15;
    assign token_in_vec_15[2] = token_2_15;
    assign in_chan_dep_vld_vec_15[3] = dep_chan_vld_3_15;
    assign in_chan_dep_data_vec_15[139 : 105] = dep_chan_data_3_15;
    assign token_in_vec_15[3] = token_3_15;
    assign in_chan_dep_vld_vec_15[4] = dep_chan_vld_4_15;
    assign in_chan_dep_data_vec_15[174 : 140] = dep_chan_data_4_15;
    assign token_in_vec_15[4] = token_4_15;
    assign in_chan_dep_vld_vec_15[5] = dep_chan_vld_5_15;
    assign in_chan_dep_data_vec_15[209 : 175] = dep_chan_data_5_15;
    assign token_in_vec_15[5] = token_5_15;
    assign in_chan_dep_vld_vec_15[6] = dep_chan_vld_6_15;
    assign in_chan_dep_data_vec_15[244 : 210] = dep_chan_data_6_15;
    assign token_in_vec_15[6] = token_6_15;
    assign in_chan_dep_vld_vec_15[7] = dep_chan_vld_7_15;
    assign in_chan_dep_data_vec_15[279 : 245] = dep_chan_data_7_15;
    assign token_in_vec_15[7] = token_7_15;
    assign in_chan_dep_vld_vec_15[8] = dep_chan_vld_8_15;
    assign in_chan_dep_data_vec_15[314 : 280] = dep_chan_data_8_15;
    assign token_in_vec_15[8] = token_8_15;
    assign in_chan_dep_vld_vec_15[9] = dep_chan_vld_9_15;
    assign in_chan_dep_data_vec_15[349 : 315] = dep_chan_data_9_15;
    assign token_in_vec_15[9] = token_9_15;
    assign in_chan_dep_vld_vec_15[10] = dep_chan_vld_10_15;
    assign in_chan_dep_data_vec_15[384 : 350] = dep_chan_data_10_15;
    assign token_in_vec_15[10] = token_10_15;
    assign in_chan_dep_vld_vec_15[11] = dep_chan_vld_11_15;
    assign in_chan_dep_data_vec_15[419 : 385] = dep_chan_data_11_15;
    assign token_in_vec_15[11] = token_11_15;
    assign in_chan_dep_vld_vec_15[12] = dep_chan_vld_12_15;
    assign in_chan_dep_data_vec_15[454 : 420] = dep_chan_data_12_15;
    assign token_in_vec_15[12] = token_12_15;
    assign in_chan_dep_vld_vec_15[13] = dep_chan_vld_13_15;
    assign in_chan_dep_data_vec_15[489 : 455] = dep_chan_data_13_15;
    assign token_in_vec_15[13] = token_13_15;
    assign in_chan_dep_vld_vec_15[14] = dep_chan_vld_14_15;
    assign in_chan_dep_data_vec_15[524 : 490] = dep_chan_data_14_15;
    assign token_in_vec_15[14] = token_14_15;
    assign in_chan_dep_vld_vec_15[15] = dep_chan_vld_16_15;
    assign in_chan_dep_data_vec_15[559 : 525] = dep_chan_data_16_15;
    assign token_in_vec_15[15] = token_16_15;
    assign in_chan_dep_vld_vec_15[16] = dep_chan_vld_17_15;
    assign in_chan_dep_data_vec_15[594 : 560] = dep_chan_data_17_15;
    assign token_in_vec_15[16] = token_17_15;
    assign in_chan_dep_vld_vec_15[17] = dep_chan_vld_18_15;
    assign in_chan_dep_data_vec_15[629 : 595] = dep_chan_data_18_15;
    assign token_in_vec_15[17] = token_18_15;
    assign in_chan_dep_vld_vec_15[18] = dep_chan_vld_31_15;
    assign in_chan_dep_data_vec_15[664 : 630] = dep_chan_data_31_15;
    assign token_in_vec_15[18] = token_31_15;
    assign dep_chan_vld_15_0 = out_chan_dep_vld_vec_15[0];
    assign dep_chan_data_15_0 = out_chan_dep_data_15;
    assign token_15_0 = token_out_vec_15[0];
    assign dep_chan_vld_15_2 = out_chan_dep_vld_vec_15[1];
    assign dep_chan_data_15_2 = out_chan_dep_data_15;
    assign token_15_2 = token_out_vec_15[1];
    assign dep_chan_vld_15_31 = out_chan_dep_vld_vec_15[2];
    assign dep_chan_data_15_31 = out_chan_dep_data_15;
    assign token_15_31 = token_out_vec_15[2];
    assign dep_chan_vld_15_1 = out_chan_dep_vld_vec_15[3];
    assign dep_chan_data_15_1 = out_chan_dep_data_15;
    assign token_15_1 = token_out_vec_15[3];
    assign dep_chan_vld_15_3 = out_chan_dep_vld_vec_15[4];
    assign dep_chan_data_15_3 = out_chan_dep_data_15;
    assign token_15_3 = token_out_vec_15[4];
    assign dep_chan_vld_15_4 = out_chan_dep_vld_vec_15[5];
    assign dep_chan_data_15_4 = out_chan_dep_data_15;
    assign token_15_4 = token_out_vec_15[5];
    assign dep_chan_vld_15_5 = out_chan_dep_vld_vec_15[6];
    assign dep_chan_data_15_5 = out_chan_dep_data_15;
    assign token_15_5 = token_out_vec_15[6];
    assign dep_chan_vld_15_6 = out_chan_dep_vld_vec_15[7];
    assign dep_chan_data_15_6 = out_chan_dep_data_15;
    assign token_15_6 = token_out_vec_15[7];
    assign dep_chan_vld_15_7 = out_chan_dep_vld_vec_15[8];
    assign dep_chan_data_15_7 = out_chan_dep_data_15;
    assign token_15_7 = token_out_vec_15[8];
    assign dep_chan_vld_15_8 = out_chan_dep_vld_vec_15[9];
    assign dep_chan_data_15_8 = out_chan_dep_data_15;
    assign token_15_8 = token_out_vec_15[9];
    assign dep_chan_vld_15_9 = out_chan_dep_vld_vec_15[10];
    assign dep_chan_data_15_9 = out_chan_dep_data_15;
    assign token_15_9 = token_out_vec_15[10];
    assign dep_chan_vld_15_10 = out_chan_dep_vld_vec_15[11];
    assign dep_chan_data_15_10 = out_chan_dep_data_15;
    assign token_15_10 = token_out_vec_15[11];
    assign dep_chan_vld_15_11 = out_chan_dep_vld_vec_15[12];
    assign dep_chan_data_15_11 = out_chan_dep_data_15;
    assign token_15_11 = token_out_vec_15[12];
    assign dep_chan_vld_15_12 = out_chan_dep_vld_vec_15[13];
    assign dep_chan_data_15_12 = out_chan_dep_data_15;
    assign token_15_12 = token_out_vec_15[13];
    assign dep_chan_vld_15_13 = out_chan_dep_vld_vec_15[14];
    assign dep_chan_data_15_13 = out_chan_dep_data_15;
    assign token_15_13 = token_out_vec_15[14];
    assign dep_chan_vld_15_14 = out_chan_dep_vld_vec_15[15];
    assign dep_chan_data_15_14 = out_chan_dep_data_15;
    assign token_15_14 = token_out_vec_15[15];
    assign dep_chan_vld_15_16 = out_chan_dep_vld_vec_15[16];
    assign dep_chan_data_15_16 = out_chan_dep_data_15;
    assign token_15_16 = token_out_vec_15[16];
    assign dep_chan_vld_15_17 = out_chan_dep_vld_vec_15[17];
    assign dep_chan_data_15_17 = out_chan_dep_data_15;
    assign token_15_17 = token_out_vec_15[17];
    assign dep_chan_vld_15_18 = out_chan_dep_vld_vec_15[18];
    assign dep_chan_data_15_18 = out_chan_dep_data_15;
    assign token_15_18 = token_out_vec_15[18];

    // Process: load_value45_U0
    kernel_pr_hls_deadlock_detect_unit #(35, 16, 19, 19) kernel_pr_hls_deadlock_detect_unit_16 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_16),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_16),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_16),
        .token_in_vec(token_in_vec_16),
        .dl_detect_in(dl_detect_out),
        .origin(origin[16]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_16),
        .out_chan_dep_data(out_chan_dep_data_16),
        .token_out_vec(token_out_vec_16),
        .dl_detect_out(dl_in_vec[16]));

    assign proc_16_data_FIFO_blk[0] = 1'b0 | (~load_value45_U0.value_r_blk_n);
    assign proc_16_data_PIPO_blk[0] = 1'b0;
    assign proc_16_start_FIFO_blk[0] = 1'b0;
    assign proc_16_TLF_FIFO_blk[0] = 1'b0;
    assign proc_16_input_sync_blk[0] = 1'b0 | (ap_sync_load_value45_U0_ap_ready & load_value45_U0.ap_idle & ~ap_sync_kernel_pr_entry98_U0_ap_ready);
    assign proc_16_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_16[0] = dl_detect_out ? proc_dep_vld_vec_16_reg[0] : (proc_16_data_FIFO_blk[0] | proc_16_data_PIPO_blk[0] | proc_16_start_FIFO_blk[0] | proc_16_TLF_FIFO_blk[0] | proc_16_input_sync_blk[0] | proc_16_output_sync_blk[0]);
    assign proc_16_data_FIFO_blk[1] = 1'b0 | (~load_value45_U0.bipedge_size_blk_n) | (~load_value45_U0.bipedge_stream_V_V13_blk_n);
    assign proc_16_data_PIPO_blk[1] = 1'b0;
    assign proc_16_start_FIFO_blk[1] = 1'b0;
    assign proc_16_TLF_FIFO_blk[1] = 1'b0;
    assign proc_16_input_sync_blk[1] = 1'b0 | (ap_sync_load_value45_U0_ap_ready & load_value45_U0.ap_idle & ~ap_sync_load_bipedge31_U0_ap_ready);
    assign proc_16_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_16[1] = dl_detect_out ? proc_dep_vld_vec_16_reg[1] : (proc_16_data_FIFO_blk[1] | proc_16_data_PIPO_blk[1] | proc_16_start_FIFO_blk[1] | proc_16_TLF_FIFO_blk[1] | proc_16_input_sync_blk[1] | proc_16_output_sync_blk[1]);
    assign proc_16_data_FIFO_blk[2] = 1'b0 | (~load_value45_U0.value_stream_V_V28_blk_n);
    assign proc_16_data_PIPO_blk[2] = 1'b0;
    assign proc_16_start_FIFO_blk[2] = 1'b0;
    assign proc_16_TLF_FIFO_blk[2] = 1'b0;
    assign proc_16_input_sync_blk[2] = 1'b0;
    assign proc_16_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_16[2] = dl_detect_out ? proc_dep_vld_vec_16_reg[2] : (proc_16_data_FIFO_blk[2] | proc_16_data_PIPO_blk[2] | proc_16_start_FIFO_blk[2] | proc_16_TLF_FIFO_blk[2] | proc_16_input_sync_blk[2] | proc_16_output_sync_blk[2]);
    assign proc_16_data_FIFO_blk[3] = 1'b0;
    assign proc_16_data_PIPO_blk[3] = 1'b0;
    assign proc_16_start_FIFO_blk[3] = 1'b0;
    assign proc_16_TLF_FIFO_blk[3] = 1'b0;
    assign proc_16_input_sync_blk[3] = 1'b0 | (ap_sync_load_value45_U0_ap_ready & load_value45_U0.ap_idle & ~ap_sync_load_bipedge30_U0_ap_ready);
    assign proc_16_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_16[3] = dl_detect_out ? proc_dep_vld_vec_16_reg[3] : (proc_16_data_FIFO_blk[3] | proc_16_data_PIPO_blk[3] | proc_16_start_FIFO_blk[3] | proc_16_TLF_FIFO_blk[3] | proc_16_input_sync_blk[3] | proc_16_output_sync_blk[3]);
    assign proc_16_data_FIFO_blk[4] = 1'b0;
    assign proc_16_data_PIPO_blk[4] = 1'b0;
    assign proc_16_start_FIFO_blk[4] = 1'b0;
    assign proc_16_TLF_FIFO_blk[4] = 1'b0;
    assign proc_16_input_sync_blk[4] = 1'b0 | (ap_sync_load_value45_U0_ap_ready & load_value45_U0.ap_idle & ~ap_sync_load_value32_U0_ap_ready);
    assign proc_16_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_16[4] = dl_detect_out ? proc_dep_vld_vec_16_reg[4] : (proc_16_data_FIFO_blk[4] | proc_16_data_PIPO_blk[4] | proc_16_start_FIFO_blk[4] | proc_16_TLF_FIFO_blk[4] | proc_16_input_sync_blk[4] | proc_16_output_sync_blk[4]);
    assign proc_16_data_FIFO_blk[5] = 1'b0;
    assign proc_16_data_PIPO_blk[5] = 1'b0;
    assign proc_16_start_FIFO_blk[5] = 1'b0;
    assign proc_16_TLF_FIFO_blk[5] = 1'b0;
    assign proc_16_input_sync_blk[5] = 1'b0 | (ap_sync_load_value45_U0_ap_ready & load_value45_U0.ap_idle & ~ap_sync_load_value33_U0_ap_ready);
    assign proc_16_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_16[5] = dl_detect_out ? proc_dep_vld_vec_16_reg[5] : (proc_16_data_FIFO_blk[5] | proc_16_data_PIPO_blk[5] | proc_16_start_FIFO_blk[5] | proc_16_TLF_FIFO_blk[5] | proc_16_input_sync_blk[5] | proc_16_output_sync_blk[5]);
    assign proc_16_data_FIFO_blk[6] = 1'b0;
    assign proc_16_data_PIPO_blk[6] = 1'b0;
    assign proc_16_start_FIFO_blk[6] = 1'b0;
    assign proc_16_TLF_FIFO_blk[6] = 1'b0;
    assign proc_16_input_sync_blk[6] = 1'b0 | (ap_sync_load_value45_U0_ap_ready & load_value45_U0.ap_idle & ~ap_sync_load_value34_U0_ap_ready);
    assign proc_16_output_sync_blk[6] = 1'b0;
    assign proc_dep_vld_vec_16[6] = dl_detect_out ? proc_dep_vld_vec_16_reg[6] : (proc_16_data_FIFO_blk[6] | proc_16_data_PIPO_blk[6] | proc_16_start_FIFO_blk[6] | proc_16_TLF_FIFO_blk[6] | proc_16_input_sync_blk[6] | proc_16_output_sync_blk[6]);
    assign proc_16_data_FIFO_blk[7] = 1'b0;
    assign proc_16_data_PIPO_blk[7] = 1'b0;
    assign proc_16_start_FIFO_blk[7] = 1'b0;
    assign proc_16_TLF_FIFO_blk[7] = 1'b0;
    assign proc_16_input_sync_blk[7] = 1'b0 | (ap_sync_load_value45_U0_ap_ready & load_value45_U0.ap_idle & ~ap_sync_load_value35_U0_ap_ready);
    assign proc_16_output_sync_blk[7] = 1'b0;
    assign proc_dep_vld_vec_16[7] = dl_detect_out ? proc_dep_vld_vec_16_reg[7] : (proc_16_data_FIFO_blk[7] | proc_16_data_PIPO_blk[7] | proc_16_start_FIFO_blk[7] | proc_16_TLF_FIFO_blk[7] | proc_16_input_sync_blk[7] | proc_16_output_sync_blk[7]);
    assign proc_16_data_FIFO_blk[8] = 1'b0;
    assign proc_16_data_PIPO_blk[8] = 1'b0;
    assign proc_16_start_FIFO_blk[8] = 1'b0;
    assign proc_16_TLF_FIFO_blk[8] = 1'b0;
    assign proc_16_input_sync_blk[8] = 1'b0 | (ap_sync_load_value45_U0_ap_ready & load_value45_U0.ap_idle & ~ap_sync_load_value36_U0_ap_ready);
    assign proc_16_output_sync_blk[8] = 1'b0;
    assign proc_dep_vld_vec_16[8] = dl_detect_out ? proc_dep_vld_vec_16_reg[8] : (proc_16_data_FIFO_blk[8] | proc_16_data_PIPO_blk[8] | proc_16_start_FIFO_blk[8] | proc_16_TLF_FIFO_blk[8] | proc_16_input_sync_blk[8] | proc_16_output_sync_blk[8]);
    assign proc_16_data_FIFO_blk[9] = 1'b0;
    assign proc_16_data_PIPO_blk[9] = 1'b0;
    assign proc_16_start_FIFO_blk[9] = 1'b0;
    assign proc_16_TLF_FIFO_blk[9] = 1'b0;
    assign proc_16_input_sync_blk[9] = 1'b0 | (ap_sync_load_value45_U0_ap_ready & load_value45_U0.ap_idle & ~ap_sync_load_value37_U0_ap_ready);
    assign proc_16_output_sync_blk[9] = 1'b0;
    assign proc_dep_vld_vec_16[9] = dl_detect_out ? proc_dep_vld_vec_16_reg[9] : (proc_16_data_FIFO_blk[9] | proc_16_data_PIPO_blk[9] | proc_16_start_FIFO_blk[9] | proc_16_TLF_FIFO_blk[9] | proc_16_input_sync_blk[9] | proc_16_output_sync_blk[9]);
    assign proc_16_data_FIFO_blk[10] = 1'b0;
    assign proc_16_data_PIPO_blk[10] = 1'b0;
    assign proc_16_start_FIFO_blk[10] = 1'b0;
    assign proc_16_TLF_FIFO_blk[10] = 1'b0;
    assign proc_16_input_sync_blk[10] = 1'b0 | (ap_sync_load_value45_U0_ap_ready & load_value45_U0.ap_idle & ~ap_sync_load_value38_U0_ap_ready);
    assign proc_16_output_sync_blk[10] = 1'b0;
    assign proc_dep_vld_vec_16[10] = dl_detect_out ? proc_dep_vld_vec_16_reg[10] : (proc_16_data_FIFO_blk[10] | proc_16_data_PIPO_blk[10] | proc_16_start_FIFO_blk[10] | proc_16_TLF_FIFO_blk[10] | proc_16_input_sync_blk[10] | proc_16_output_sync_blk[10]);
    assign proc_16_data_FIFO_blk[11] = 1'b0;
    assign proc_16_data_PIPO_blk[11] = 1'b0;
    assign proc_16_start_FIFO_blk[11] = 1'b0;
    assign proc_16_TLF_FIFO_blk[11] = 1'b0;
    assign proc_16_input_sync_blk[11] = 1'b0 | (ap_sync_load_value45_U0_ap_ready & load_value45_U0.ap_idle & ~ap_sync_load_value39_U0_ap_ready);
    assign proc_16_output_sync_blk[11] = 1'b0;
    assign proc_dep_vld_vec_16[11] = dl_detect_out ? proc_dep_vld_vec_16_reg[11] : (proc_16_data_FIFO_blk[11] | proc_16_data_PIPO_blk[11] | proc_16_start_FIFO_blk[11] | proc_16_TLF_FIFO_blk[11] | proc_16_input_sync_blk[11] | proc_16_output_sync_blk[11]);
    assign proc_16_data_FIFO_blk[12] = 1'b0;
    assign proc_16_data_PIPO_blk[12] = 1'b0;
    assign proc_16_start_FIFO_blk[12] = 1'b0;
    assign proc_16_TLF_FIFO_blk[12] = 1'b0;
    assign proc_16_input_sync_blk[12] = 1'b0 | (ap_sync_load_value45_U0_ap_ready & load_value45_U0.ap_idle & ~ap_sync_load_value40_U0_ap_ready);
    assign proc_16_output_sync_blk[12] = 1'b0;
    assign proc_dep_vld_vec_16[12] = dl_detect_out ? proc_dep_vld_vec_16_reg[12] : (proc_16_data_FIFO_blk[12] | proc_16_data_PIPO_blk[12] | proc_16_start_FIFO_blk[12] | proc_16_TLF_FIFO_blk[12] | proc_16_input_sync_blk[12] | proc_16_output_sync_blk[12]);
    assign proc_16_data_FIFO_blk[13] = 1'b0;
    assign proc_16_data_PIPO_blk[13] = 1'b0;
    assign proc_16_start_FIFO_blk[13] = 1'b0;
    assign proc_16_TLF_FIFO_blk[13] = 1'b0;
    assign proc_16_input_sync_blk[13] = 1'b0 | (ap_sync_load_value45_U0_ap_ready & load_value45_U0.ap_idle & ~ap_sync_load_value41_U0_ap_ready);
    assign proc_16_output_sync_blk[13] = 1'b0;
    assign proc_dep_vld_vec_16[13] = dl_detect_out ? proc_dep_vld_vec_16_reg[13] : (proc_16_data_FIFO_blk[13] | proc_16_data_PIPO_blk[13] | proc_16_start_FIFO_blk[13] | proc_16_TLF_FIFO_blk[13] | proc_16_input_sync_blk[13] | proc_16_output_sync_blk[13]);
    assign proc_16_data_FIFO_blk[14] = 1'b0;
    assign proc_16_data_PIPO_blk[14] = 1'b0;
    assign proc_16_start_FIFO_blk[14] = 1'b0;
    assign proc_16_TLF_FIFO_blk[14] = 1'b0;
    assign proc_16_input_sync_blk[14] = 1'b0 | (ap_sync_load_value45_U0_ap_ready & load_value45_U0.ap_idle & ~ap_sync_load_value42_U0_ap_ready);
    assign proc_16_output_sync_blk[14] = 1'b0;
    assign proc_dep_vld_vec_16[14] = dl_detect_out ? proc_dep_vld_vec_16_reg[14] : (proc_16_data_FIFO_blk[14] | proc_16_data_PIPO_blk[14] | proc_16_start_FIFO_blk[14] | proc_16_TLF_FIFO_blk[14] | proc_16_input_sync_blk[14] | proc_16_output_sync_blk[14]);
    assign proc_16_data_FIFO_blk[15] = 1'b0;
    assign proc_16_data_PIPO_blk[15] = 1'b0;
    assign proc_16_start_FIFO_blk[15] = 1'b0;
    assign proc_16_TLF_FIFO_blk[15] = 1'b0;
    assign proc_16_input_sync_blk[15] = 1'b0 | (ap_sync_load_value45_U0_ap_ready & load_value45_U0.ap_idle & ~ap_sync_load_value43_U0_ap_ready);
    assign proc_16_output_sync_blk[15] = 1'b0;
    assign proc_dep_vld_vec_16[15] = dl_detect_out ? proc_dep_vld_vec_16_reg[15] : (proc_16_data_FIFO_blk[15] | proc_16_data_PIPO_blk[15] | proc_16_start_FIFO_blk[15] | proc_16_TLF_FIFO_blk[15] | proc_16_input_sync_blk[15] | proc_16_output_sync_blk[15]);
    assign proc_16_data_FIFO_blk[16] = 1'b0;
    assign proc_16_data_PIPO_blk[16] = 1'b0;
    assign proc_16_start_FIFO_blk[16] = 1'b0;
    assign proc_16_TLF_FIFO_blk[16] = 1'b0;
    assign proc_16_input_sync_blk[16] = 1'b0 | (ap_sync_load_value45_U0_ap_ready & load_value45_U0.ap_idle & ~ap_sync_load_value44_U0_ap_ready);
    assign proc_16_output_sync_blk[16] = 1'b0;
    assign proc_dep_vld_vec_16[16] = dl_detect_out ? proc_dep_vld_vec_16_reg[16] : (proc_16_data_FIFO_blk[16] | proc_16_data_PIPO_blk[16] | proc_16_start_FIFO_blk[16] | proc_16_TLF_FIFO_blk[16] | proc_16_input_sync_blk[16] | proc_16_output_sync_blk[16]);
    assign proc_16_data_FIFO_blk[17] = 1'b0;
    assign proc_16_data_PIPO_blk[17] = 1'b0;
    assign proc_16_start_FIFO_blk[17] = 1'b0;
    assign proc_16_TLF_FIFO_blk[17] = 1'b0;
    assign proc_16_input_sync_blk[17] = 1'b0 | (ap_sync_load_value45_U0_ap_ready & load_value45_U0.ap_idle & ~ap_sync_load_value46_U0_ap_ready);
    assign proc_16_output_sync_blk[17] = 1'b0;
    assign proc_dep_vld_vec_16[17] = dl_detect_out ? proc_dep_vld_vec_16_reg[17] : (proc_16_data_FIFO_blk[17] | proc_16_data_PIPO_blk[17] | proc_16_start_FIFO_blk[17] | proc_16_TLF_FIFO_blk[17] | proc_16_input_sync_blk[17] | proc_16_output_sync_blk[17]);
    assign proc_16_data_FIFO_blk[18] = 1'b0;
    assign proc_16_data_PIPO_blk[18] = 1'b0;
    assign proc_16_start_FIFO_blk[18] = 1'b0;
    assign proc_16_TLF_FIFO_blk[18] = 1'b0;
    assign proc_16_input_sync_blk[18] = 1'b0 | (ap_sync_load_value45_U0_ap_ready & load_value45_U0.ap_idle & ~ap_sync_load_value47_U0_ap_ready);
    assign proc_16_output_sync_blk[18] = 1'b0;
    assign proc_dep_vld_vec_16[18] = dl_detect_out ? proc_dep_vld_vec_16_reg[18] : (proc_16_data_FIFO_blk[18] | proc_16_data_PIPO_blk[18] | proc_16_start_FIFO_blk[18] | proc_16_TLF_FIFO_blk[18] | proc_16_input_sync_blk[18] | proc_16_output_sync_blk[18]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_16_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_16_reg <= proc_dep_vld_vec_16;
        end
    end
    assign in_chan_dep_vld_vec_16[0] = dep_chan_vld_0_16;
    assign in_chan_dep_data_vec_16[34 : 0] = dep_chan_data_0_16;
    assign token_in_vec_16[0] = token_0_16;
    assign in_chan_dep_vld_vec_16[1] = dep_chan_vld_1_16;
    assign in_chan_dep_data_vec_16[69 : 35] = dep_chan_data_1_16;
    assign token_in_vec_16[1] = token_1_16;
    assign in_chan_dep_vld_vec_16[2] = dep_chan_vld_2_16;
    assign in_chan_dep_data_vec_16[104 : 70] = dep_chan_data_2_16;
    assign token_in_vec_16[2] = token_2_16;
    assign in_chan_dep_vld_vec_16[3] = dep_chan_vld_3_16;
    assign in_chan_dep_data_vec_16[139 : 105] = dep_chan_data_3_16;
    assign token_in_vec_16[3] = token_3_16;
    assign in_chan_dep_vld_vec_16[4] = dep_chan_vld_4_16;
    assign in_chan_dep_data_vec_16[174 : 140] = dep_chan_data_4_16;
    assign token_in_vec_16[4] = token_4_16;
    assign in_chan_dep_vld_vec_16[5] = dep_chan_vld_5_16;
    assign in_chan_dep_data_vec_16[209 : 175] = dep_chan_data_5_16;
    assign token_in_vec_16[5] = token_5_16;
    assign in_chan_dep_vld_vec_16[6] = dep_chan_vld_6_16;
    assign in_chan_dep_data_vec_16[244 : 210] = dep_chan_data_6_16;
    assign token_in_vec_16[6] = token_6_16;
    assign in_chan_dep_vld_vec_16[7] = dep_chan_vld_7_16;
    assign in_chan_dep_data_vec_16[279 : 245] = dep_chan_data_7_16;
    assign token_in_vec_16[7] = token_7_16;
    assign in_chan_dep_vld_vec_16[8] = dep_chan_vld_8_16;
    assign in_chan_dep_data_vec_16[314 : 280] = dep_chan_data_8_16;
    assign token_in_vec_16[8] = token_8_16;
    assign in_chan_dep_vld_vec_16[9] = dep_chan_vld_9_16;
    assign in_chan_dep_data_vec_16[349 : 315] = dep_chan_data_9_16;
    assign token_in_vec_16[9] = token_9_16;
    assign in_chan_dep_vld_vec_16[10] = dep_chan_vld_10_16;
    assign in_chan_dep_data_vec_16[384 : 350] = dep_chan_data_10_16;
    assign token_in_vec_16[10] = token_10_16;
    assign in_chan_dep_vld_vec_16[11] = dep_chan_vld_11_16;
    assign in_chan_dep_data_vec_16[419 : 385] = dep_chan_data_11_16;
    assign token_in_vec_16[11] = token_11_16;
    assign in_chan_dep_vld_vec_16[12] = dep_chan_vld_12_16;
    assign in_chan_dep_data_vec_16[454 : 420] = dep_chan_data_12_16;
    assign token_in_vec_16[12] = token_12_16;
    assign in_chan_dep_vld_vec_16[13] = dep_chan_vld_13_16;
    assign in_chan_dep_data_vec_16[489 : 455] = dep_chan_data_13_16;
    assign token_in_vec_16[13] = token_13_16;
    assign in_chan_dep_vld_vec_16[14] = dep_chan_vld_14_16;
    assign in_chan_dep_data_vec_16[524 : 490] = dep_chan_data_14_16;
    assign token_in_vec_16[14] = token_14_16;
    assign in_chan_dep_vld_vec_16[15] = dep_chan_vld_15_16;
    assign in_chan_dep_data_vec_16[559 : 525] = dep_chan_data_15_16;
    assign token_in_vec_16[15] = token_15_16;
    assign in_chan_dep_vld_vec_16[16] = dep_chan_vld_17_16;
    assign in_chan_dep_data_vec_16[594 : 560] = dep_chan_data_17_16;
    assign token_in_vec_16[16] = token_17_16;
    assign in_chan_dep_vld_vec_16[17] = dep_chan_vld_18_16;
    assign in_chan_dep_data_vec_16[629 : 595] = dep_chan_data_18_16;
    assign token_in_vec_16[17] = token_18_16;
    assign in_chan_dep_vld_vec_16[18] = dep_chan_vld_32_16;
    assign in_chan_dep_data_vec_16[664 : 630] = dep_chan_data_32_16;
    assign token_in_vec_16[18] = token_32_16;
    assign dep_chan_vld_16_0 = out_chan_dep_vld_vec_16[0];
    assign dep_chan_data_16_0 = out_chan_dep_data_16;
    assign token_16_0 = token_out_vec_16[0];
    assign dep_chan_vld_16_2 = out_chan_dep_vld_vec_16[1];
    assign dep_chan_data_16_2 = out_chan_dep_data_16;
    assign token_16_2 = token_out_vec_16[1];
    assign dep_chan_vld_16_32 = out_chan_dep_vld_vec_16[2];
    assign dep_chan_data_16_32 = out_chan_dep_data_16;
    assign token_16_32 = token_out_vec_16[2];
    assign dep_chan_vld_16_1 = out_chan_dep_vld_vec_16[3];
    assign dep_chan_data_16_1 = out_chan_dep_data_16;
    assign token_16_1 = token_out_vec_16[3];
    assign dep_chan_vld_16_3 = out_chan_dep_vld_vec_16[4];
    assign dep_chan_data_16_3 = out_chan_dep_data_16;
    assign token_16_3 = token_out_vec_16[4];
    assign dep_chan_vld_16_4 = out_chan_dep_vld_vec_16[5];
    assign dep_chan_data_16_4 = out_chan_dep_data_16;
    assign token_16_4 = token_out_vec_16[5];
    assign dep_chan_vld_16_5 = out_chan_dep_vld_vec_16[6];
    assign dep_chan_data_16_5 = out_chan_dep_data_16;
    assign token_16_5 = token_out_vec_16[6];
    assign dep_chan_vld_16_6 = out_chan_dep_vld_vec_16[7];
    assign dep_chan_data_16_6 = out_chan_dep_data_16;
    assign token_16_6 = token_out_vec_16[7];
    assign dep_chan_vld_16_7 = out_chan_dep_vld_vec_16[8];
    assign dep_chan_data_16_7 = out_chan_dep_data_16;
    assign token_16_7 = token_out_vec_16[8];
    assign dep_chan_vld_16_8 = out_chan_dep_vld_vec_16[9];
    assign dep_chan_data_16_8 = out_chan_dep_data_16;
    assign token_16_8 = token_out_vec_16[9];
    assign dep_chan_vld_16_9 = out_chan_dep_vld_vec_16[10];
    assign dep_chan_data_16_9 = out_chan_dep_data_16;
    assign token_16_9 = token_out_vec_16[10];
    assign dep_chan_vld_16_10 = out_chan_dep_vld_vec_16[11];
    assign dep_chan_data_16_10 = out_chan_dep_data_16;
    assign token_16_10 = token_out_vec_16[11];
    assign dep_chan_vld_16_11 = out_chan_dep_vld_vec_16[12];
    assign dep_chan_data_16_11 = out_chan_dep_data_16;
    assign token_16_11 = token_out_vec_16[12];
    assign dep_chan_vld_16_12 = out_chan_dep_vld_vec_16[13];
    assign dep_chan_data_16_12 = out_chan_dep_data_16;
    assign token_16_12 = token_out_vec_16[13];
    assign dep_chan_vld_16_13 = out_chan_dep_vld_vec_16[14];
    assign dep_chan_data_16_13 = out_chan_dep_data_16;
    assign token_16_13 = token_out_vec_16[14];
    assign dep_chan_vld_16_14 = out_chan_dep_vld_vec_16[15];
    assign dep_chan_data_16_14 = out_chan_dep_data_16;
    assign token_16_14 = token_out_vec_16[15];
    assign dep_chan_vld_16_15 = out_chan_dep_vld_vec_16[16];
    assign dep_chan_data_16_15 = out_chan_dep_data_16;
    assign token_16_15 = token_out_vec_16[16];
    assign dep_chan_vld_16_17 = out_chan_dep_vld_vec_16[17];
    assign dep_chan_data_16_17 = out_chan_dep_data_16;
    assign token_16_17 = token_out_vec_16[17];
    assign dep_chan_vld_16_18 = out_chan_dep_vld_vec_16[18];
    assign dep_chan_data_16_18 = out_chan_dep_data_16;
    assign token_16_18 = token_out_vec_16[18];

    // Process: load_value46_U0
    kernel_pr_hls_deadlock_detect_unit #(35, 17, 19, 19) kernel_pr_hls_deadlock_detect_unit_17 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_17),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_17),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_17),
        .token_in_vec(token_in_vec_17),
        .dl_detect_in(dl_detect_out),
        .origin(origin[17]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_17),
        .out_chan_dep_data(out_chan_dep_data_17),
        .token_out_vec(token_out_vec_17),
        .dl_detect_out(dl_in_vec[17]));

    assign proc_17_data_FIFO_blk[0] = 1'b0 | (~load_value46_U0.value_r_blk_n);
    assign proc_17_data_PIPO_blk[0] = 1'b0;
    assign proc_17_start_FIFO_blk[0] = 1'b0;
    assign proc_17_TLF_FIFO_blk[0] = 1'b0;
    assign proc_17_input_sync_blk[0] = 1'b0 | (ap_sync_load_value46_U0_ap_ready & load_value46_U0.ap_idle & ~ap_sync_kernel_pr_entry98_U0_ap_ready);
    assign proc_17_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_17[0] = dl_detect_out ? proc_dep_vld_vec_17_reg[0] : (proc_17_data_FIFO_blk[0] | proc_17_data_PIPO_blk[0] | proc_17_start_FIFO_blk[0] | proc_17_TLF_FIFO_blk[0] | proc_17_input_sync_blk[0] | proc_17_output_sync_blk[0]);
    assign proc_17_data_FIFO_blk[1] = 1'b0 | (~load_value46_U0.bipedge_size_blk_n) | (~load_value46_U0.bipedge_stream_V_V14_blk_n);
    assign proc_17_data_PIPO_blk[1] = 1'b0;
    assign proc_17_start_FIFO_blk[1] = 1'b0;
    assign proc_17_TLF_FIFO_blk[1] = 1'b0;
    assign proc_17_input_sync_blk[1] = 1'b0 | (ap_sync_load_value46_U0_ap_ready & load_value46_U0.ap_idle & ~ap_sync_load_bipedge31_U0_ap_ready);
    assign proc_17_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_17[1] = dl_detect_out ? proc_dep_vld_vec_17_reg[1] : (proc_17_data_FIFO_blk[1] | proc_17_data_PIPO_blk[1] | proc_17_start_FIFO_blk[1] | proc_17_TLF_FIFO_blk[1] | proc_17_input_sync_blk[1] | proc_17_output_sync_blk[1]);
    assign proc_17_data_FIFO_blk[2] = 1'b0 | (~load_value46_U0.value_stream_V_V29_blk_n);
    assign proc_17_data_PIPO_blk[2] = 1'b0;
    assign proc_17_start_FIFO_blk[2] = 1'b0;
    assign proc_17_TLF_FIFO_blk[2] = 1'b0;
    assign proc_17_input_sync_blk[2] = 1'b0;
    assign proc_17_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_17[2] = dl_detect_out ? proc_dep_vld_vec_17_reg[2] : (proc_17_data_FIFO_blk[2] | proc_17_data_PIPO_blk[2] | proc_17_start_FIFO_blk[2] | proc_17_TLF_FIFO_blk[2] | proc_17_input_sync_blk[2] | proc_17_output_sync_blk[2]);
    assign proc_17_data_FIFO_blk[3] = 1'b0;
    assign proc_17_data_PIPO_blk[3] = 1'b0;
    assign proc_17_start_FIFO_blk[3] = 1'b0;
    assign proc_17_TLF_FIFO_blk[3] = 1'b0;
    assign proc_17_input_sync_blk[3] = 1'b0 | (ap_sync_load_value46_U0_ap_ready & load_value46_U0.ap_idle & ~ap_sync_load_bipedge30_U0_ap_ready);
    assign proc_17_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_17[3] = dl_detect_out ? proc_dep_vld_vec_17_reg[3] : (proc_17_data_FIFO_blk[3] | proc_17_data_PIPO_blk[3] | proc_17_start_FIFO_blk[3] | proc_17_TLF_FIFO_blk[3] | proc_17_input_sync_blk[3] | proc_17_output_sync_blk[3]);
    assign proc_17_data_FIFO_blk[4] = 1'b0;
    assign proc_17_data_PIPO_blk[4] = 1'b0;
    assign proc_17_start_FIFO_blk[4] = 1'b0;
    assign proc_17_TLF_FIFO_blk[4] = 1'b0;
    assign proc_17_input_sync_blk[4] = 1'b0 | (ap_sync_load_value46_U0_ap_ready & load_value46_U0.ap_idle & ~ap_sync_load_value32_U0_ap_ready);
    assign proc_17_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_17[4] = dl_detect_out ? proc_dep_vld_vec_17_reg[4] : (proc_17_data_FIFO_blk[4] | proc_17_data_PIPO_blk[4] | proc_17_start_FIFO_blk[4] | proc_17_TLF_FIFO_blk[4] | proc_17_input_sync_blk[4] | proc_17_output_sync_blk[4]);
    assign proc_17_data_FIFO_blk[5] = 1'b0;
    assign proc_17_data_PIPO_blk[5] = 1'b0;
    assign proc_17_start_FIFO_blk[5] = 1'b0;
    assign proc_17_TLF_FIFO_blk[5] = 1'b0;
    assign proc_17_input_sync_blk[5] = 1'b0 | (ap_sync_load_value46_U0_ap_ready & load_value46_U0.ap_idle & ~ap_sync_load_value33_U0_ap_ready);
    assign proc_17_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_17[5] = dl_detect_out ? proc_dep_vld_vec_17_reg[5] : (proc_17_data_FIFO_blk[5] | proc_17_data_PIPO_blk[5] | proc_17_start_FIFO_blk[5] | proc_17_TLF_FIFO_blk[5] | proc_17_input_sync_blk[5] | proc_17_output_sync_blk[5]);
    assign proc_17_data_FIFO_blk[6] = 1'b0;
    assign proc_17_data_PIPO_blk[6] = 1'b0;
    assign proc_17_start_FIFO_blk[6] = 1'b0;
    assign proc_17_TLF_FIFO_blk[6] = 1'b0;
    assign proc_17_input_sync_blk[6] = 1'b0 | (ap_sync_load_value46_U0_ap_ready & load_value46_U0.ap_idle & ~ap_sync_load_value34_U0_ap_ready);
    assign proc_17_output_sync_blk[6] = 1'b0;
    assign proc_dep_vld_vec_17[6] = dl_detect_out ? proc_dep_vld_vec_17_reg[6] : (proc_17_data_FIFO_blk[6] | proc_17_data_PIPO_blk[6] | proc_17_start_FIFO_blk[6] | proc_17_TLF_FIFO_blk[6] | proc_17_input_sync_blk[6] | proc_17_output_sync_blk[6]);
    assign proc_17_data_FIFO_blk[7] = 1'b0;
    assign proc_17_data_PIPO_blk[7] = 1'b0;
    assign proc_17_start_FIFO_blk[7] = 1'b0;
    assign proc_17_TLF_FIFO_blk[7] = 1'b0;
    assign proc_17_input_sync_blk[7] = 1'b0 | (ap_sync_load_value46_U0_ap_ready & load_value46_U0.ap_idle & ~ap_sync_load_value35_U0_ap_ready);
    assign proc_17_output_sync_blk[7] = 1'b0;
    assign proc_dep_vld_vec_17[7] = dl_detect_out ? proc_dep_vld_vec_17_reg[7] : (proc_17_data_FIFO_blk[7] | proc_17_data_PIPO_blk[7] | proc_17_start_FIFO_blk[7] | proc_17_TLF_FIFO_blk[7] | proc_17_input_sync_blk[7] | proc_17_output_sync_blk[7]);
    assign proc_17_data_FIFO_blk[8] = 1'b0;
    assign proc_17_data_PIPO_blk[8] = 1'b0;
    assign proc_17_start_FIFO_blk[8] = 1'b0;
    assign proc_17_TLF_FIFO_blk[8] = 1'b0;
    assign proc_17_input_sync_blk[8] = 1'b0 | (ap_sync_load_value46_U0_ap_ready & load_value46_U0.ap_idle & ~ap_sync_load_value36_U0_ap_ready);
    assign proc_17_output_sync_blk[8] = 1'b0;
    assign proc_dep_vld_vec_17[8] = dl_detect_out ? proc_dep_vld_vec_17_reg[8] : (proc_17_data_FIFO_blk[8] | proc_17_data_PIPO_blk[8] | proc_17_start_FIFO_blk[8] | proc_17_TLF_FIFO_blk[8] | proc_17_input_sync_blk[8] | proc_17_output_sync_blk[8]);
    assign proc_17_data_FIFO_blk[9] = 1'b0;
    assign proc_17_data_PIPO_blk[9] = 1'b0;
    assign proc_17_start_FIFO_blk[9] = 1'b0;
    assign proc_17_TLF_FIFO_blk[9] = 1'b0;
    assign proc_17_input_sync_blk[9] = 1'b0 | (ap_sync_load_value46_U0_ap_ready & load_value46_U0.ap_idle & ~ap_sync_load_value37_U0_ap_ready);
    assign proc_17_output_sync_blk[9] = 1'b0;
    assign proc_dep_vld_vec_17[9] = dl_detect_out ? proc_dep_vld_vec_17_reg[9] : (proc_17_data_FIFO_blk[9] | proc_17_data_PIPO_blk[9] | proc_17_start_FIFO_blk[9] | proc_17_TLF_FIFO_blk[9] | proc_17_input_sync_blk[9] | proc_17_output_sync_blk[9]);
    assign proc_17_data_FIFO_blk[10] = 1'b0;
    assign proc_17_data_PIPO_blk[10] = 1'b0;
    assign proc_17_start_FIFO_blk[10] = 1'b0;
    assign proc_17_TLF_FIFO_blk[10] = 1'b0;
    assign proc_17_input_sync_blk[10] = 1'b0 | (ap_sync_load_value46_U0_ap_ready & load_value46_U0.ap_idle & ~ap_sync_load_value38_U0_ap_ready);
    assign proc_17_output_sync_blk[10] = 1'b0;
    assign proc_dep_vld_vec_17[10] = dl_detect_out ? proc_dep_vld_vec_17_reg[10] : (proc_17_data_FIFO_blk[10] | proc_17_data_PIPO_blk[10] | proc_17_start_FIFO_blk[10] | proc_17_TLF_FIFO_blk[10] | proc_17_input_sync_blk[10] | proc_17_output_sync_blk[10]);
    assign proc_17_data_FIFO_blk[11] = 1'b0;
    assign proc_17_data_PIPO_blk[11] = 1'b0;
    assign proc_17_start_FIFO_blk[11] = 1'b0;
    assign proc_17_TLF_FIFO_blk[11] = 1'b0;
    assign proc_17_input_sync_blk[11] = 1'b0 | (ap_sync_load_value46_U0_ap_ready & load_value46_U0.ap_idle & ~ap_sync_load_value39_U0_ap_ready);
    assign proc_17_output_sync_blk[11] = 1'b0;
    assign proc_dep_vld_vec_17[11] = dl_detect_out ? proc_dep_vld_vec_17_reg[11] : (proc_17_data_FIFO_blk[11] | proc_17_data_PIPO_blk[11] | proc_17_start_FIFO_blk[11] | proc_17_TLF_FIFO_blk[11] | proc_17_input_sync_blk[11] | proc_17_output_sync_blk[11]);
    assign proc_17_data_FIFO_blk[12] = 1'b0;
    assign proc_17_data_PIPO_blk[12] = 1'b0;
    assign proc_17_start_FIFO_blk[12] = 1'b0;
    assign proc_17_TLF_FIFO_blk[12] = 1'b0;
    assign proc_17_input_sync_blk[12] = 1'b0 | (ap_sync_load_value46_U0_ap_ready & load_value46_U0.ap_idle & ~ap_sync_load_value40_U0_ap_ready);
    assign proc_17_output_sync_blk[12] = 1'b0;
    assign proc_dep_vld_vec_17[12] = dl_detect_out ? proc_dep_vld_vec_17_reg[12] : (proc_17_data_FIFO_blk[12] | proc_17_data_PIPO_blk[12] | proc_17_start_FIFO_blk[12] | proc_17_TLF_FIFO_blk[12] | proc_17_input_sync_blk[12] | proc_17_output_sync_blk[12]);
    assign proc_17_data_FIFO_blk[13] = 1'b0;
    assign proc_17_data_PIPO_blk[13] = 1'b0;
    assign proc_17_start_FIFO_blk[13] = 1'b0;
    assign proc_17_TLF_FIFO_blk[13] = 1'b0;
    assign proc_17_input_sync_blk[13] = 1'b0 | (ap_sync_load_value46_U0_ap_ready & load_value46_U0.ap_idle & ~ap_sync_load_value41_U0_ap_ready);
    assign proc_17_output_sync_blk[13] = 1'b0;
    assign proc_dep_vld_vec_17[13] = dl_detect_out ? proc_dep_vld_vec_17_reg[13] : (proc_17_data_FIFO_blk[13] | proc_17_data_PIPO_blk[13] | proc_17_start_FIFO_blk[13] | proc_17_TLF_FIFO_blk[13] | proc_17_input_sync_blk[13] | proc_17_output_sync_blk[13]);
    assign proc_17_data_FIFO_blk[14] = 1'b0;
    assign proc_17_data_PIPO_blk[14] = 1'b0;
    assign proc_17_start_FIFO_blk[14] = 1'b0;
    assign proc_17_TLF_FIFO_blk[14] = 1'b0;
    assign proc_17_input_sync_blk[14] = 1'b0 | (ap_sync_load_value46_U0_ap_ready & load_value46_U0.ap_idle & ~ap_sync_load_value42_U0_ap_ready);
    assign proc_17_output_sync_blk[14] = 1'b0;
    assign proc_dep_vld_vec_17[14] = dl_detect_out ? proc_dep_vld_vec_17_reg[14] : (proc_17_data_FIFO_blk[14] | proc_17_data_PIPO_blk[14] | proc_17_start_FIFO_blk[14] | proc_17_TLF_FIFO_blk[14] | proc_17_input_sync_blk[14] | proc_17_output_sync_blk[14]);
    assign proc_17_data_FIFO_blk[15] = 1'b0;
    assign proc_17_data_PIPO_blk[15] = 1'b0;
    assign proc_17_start_FIFO_blk[15] = 1'b0;
    assign proc_17_TLF_FIFO_blk[15] = 1'b0;
    assign proc_17_input_sync_blk[15] = 1'b0 | (ap_sync_load_value46_U0_ap_ready & load_value46_U0.ap_idle & ~ap_sync_load_value43_U0_ap_ready);
    assign proc_17_output_sync_blk[15] = 1'b0;
    assign proc_dep_vld_vec_17[15] = dl_detect_out ? proc_dep_vld_vec_17_reg[15] : (proc_17_data_FIFO_blk[15] | proc_17_data_PIPO_blk[15] | proc_17_start_FIFO_blk[15] | proc_17_TLF_FIFO_blk[15] | proc_17_input_sync_blk[15] | proc_17_output_sync_blk[15]);
    assign proc_17_data_FIFO_blk[16] = 1'b0;
    assign proc_17_data_PIPO_blk[16] = 1'b0;
    assign proc_17_start_FIFO_blk[16] = 1'b0;
    assign proc_17_TLF_FIFO_blk[16] = 1'b0;
    assign proc_17_input_sync_blk[16] = 1'b0 | (ap_sync_load_value46_U0_ap_ready & load_value46_U0.ap_idle & ~ap_sync_load_value44_U0_ap_ready);
    assign proc_17_output_sync_blk[16] = 1'b0;
    assign proc_dep_vld_vec_17[16] = dl_detect_out ? proc_dep_vld_vec_17_reg[16] : (proc_17_data_FIFO_blk[16] | proc_17_data_PIPO_blk[16] | proc_17_start_FIFO_blk[16] | proc_17_TLF_FIFO_blk[16] | proc_17_input_sync_blk[16] | proc_17_output_sync_blk[16]);
    assign proc_17_data_FIFO_blk[17] = 1'b0;
    assign proc_17_data_PIPO_blk[17] = 1'b0;
    assign proc_17_start_FIFO_blk[17] = 1'b0;
    assign proc_17_TLF_FIFO_blk[17] = 1'b0;
    assign proc_17_input_sync_blk[17] = 1'b0 | (ap_sync_load_value46_U0_ap_ready & load_value46_U0.ap_idle & ~ap_sync_load_value45_U0_ap_ready);
    assign proc_17_output_sync_blk[17] = 1'b0;
    assign proc_dep_vld_vec_17[17] = dl_detect_out ? proc_dep_vld_vec_17_reg[17] : (proc_17_data_FIFO_blk[17] | proc_17_data_PIPO_blk[17] | proc_17_start_FIFO_blk[17] | proc_17_TLF_FIFO_blk[17] | proc_17_input_sync_blk[17] | proc_17_output_sync_blk[17]);
    assign proc_17_data_FIFO_blk[18] = 1'b0;
    assign proc_17_data_PIPO_blk[18] = 1'b0;
    assign proc_17_start_FIFO_blk[18] = 1'b0;
    assign proc_17_TLF_FIFO_blk[18] = 1'b0;
    assign proc_17_input_sync_blk[18] = 1'b0 | (ap_sync_load_value46_U0_ap_ready & load_value46_U0.ap_idle & ~ap_sync_load_value47_U0_ap_ready);
    assign proc_17_output_sync_blk[18] = 1'b0;
    assign proc_dep_vld_vec_17[18] = dl_detect_out ? proc_dep_vld_vec_17_reg[18] : (proc_17_data_FIFO_blk[18] | proc_17_data_PIPO_blk[18] | proc_17_start_FIFO_blk[18] | proc_17_TLF_FIFO_blk[18] | proc_17_input_sync_blk[18] | proc_17_output_sync_blk[18]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_17_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_17_reg <= proc_dep_vld_vec_17;
        end
    end
    assign in_chan_dep_vld_vec_17[0] = dep_chan_vld_0_17;
    assign in_chan_dep_data_vec_17[34 : 0] = dep_chan_data_0_17;
    assign token_in_vec_17[0] = token_0_17;
    assign in_chan_dep_vld_vec_17[1] = dep_chan_vld_1_17;
    assign in_chan_dep_data_vec_17[69 : 35] = dep_chan_data_1_17;
    assign token_in_vec_17[1] = token_1_17;
    assign in_chan_dep_vld_vec_17[2] = dep_chan_vld_2_17;
    assign in_chan_dep_data_vec_17[104 : 70] = dep_chan_data_2_17;
    assign token_in_vec_17[2] = token_2_17;
    assign in_chan_dep_vld_vec_17[3] = dep_chan_vld_3_17;
    assign in_chan_dep_data_vec_17[139 : 105] = dep_chan_data_3_17;
    assign token_in_vec_17[3] = token_3_17;
    assign in_chan_dep_vld_vec_17[4] = dep_chan_vld_4_17;
    assign in_chan_dep_data_vec_17[174 : 140] = dep_chan_data_4_17;
    assign token_in_vec_17[4] = token_4_17;
    assign in_chan_dep_vld_vec_17[5] = dep_chan_vld_5_17;
    assign in_chan_dep_data_vec_17[209 : 175] = dep_chan_data_5_17;
    assign token_in_vec_17[5] = token_5_17;
    assign in_chan_dep_vld_vec_17[6] = dep_chan_vld_6_17;
    assign in_chan_dep_data_vec_17[244 : 210] = dep_chan_data_6_17;
    assign token_in_vec_17[6] = token_6_17;
    assign in_chan_dep_vld_vec_17[7] = dep_chan_vld_7_17;
    assign in_chan_dep_data_vec_17[279 : 245] = dep_chan_data_7_17;
    assign token_in_vec_17[7] = token_7_17;
    assign in_chan_dep_vld_vec_17[8] = dep_chan_vld_8_17;
    assign in_chan_dep_data_vec_17[314 : 280] = dep_chan_data_8_17;
    assign token_in_vec_17[8] = token_8_17;
    assign in_chan_dep_vld_vec_17[9] = dep_chan_vld_9_17;
    assign in_chan_dep_data_vec_17[349 : 315] = dep_chan_data_9_17;
    assign token_in_vec_17[9] = token_9_17;
    assign in_chan_dep_vld_vec_17[10] = dep_chan_vld_10_17;
    assign in_chan_dep_data_vec_17[384 : 350] = dep_chan_data_10_17;
    assign token_in_vec_17[10] = token_10_17;
    assign in_chan_dep_vld_vec_17[11] = dep_chan_vld_11_17;
    assign in_chan_dep_data_vec_17[419 : 385] = dep_chan_data_11_17;
    assign token_in_vec_17[11] = token_11_17;
    assign in_chan_dep_vld_vec_17[12] = dep_chan_vld_12_17;
    assign in_chan_dep_data_vec_17[454 : 420] = dep_chan_data_12_17;
    assign token_in_vec_17[12] = token_12_17;
    assign in_chan_dep_vld_vec_17[13] = dep_chan_vld_13_17;
    assign in_chan_dep_data_vec_17[489 : 455] = dep_chan_data_13_17;
    assign token_in_vec_17[13] = token_13_17;
    assign in_chan_dep_vld_vec_17[14] = dep_chan_vld_14_17;
    assign in_chan_dep_data_vec_17[524 : 490] = dep_chan_data_14_17;
    assign token_in_vec_17[14] = token_14_17;
    assign in_chan_dep_vld_vec_17[15] = dep_chan_vld_15_17;
    assign in_chan_dep_data_vec_17[559 : 525] = dep_chan_data_15_17;
    assign token_in_vec_17[15] = token_15_17;
    assign in_chan_dep_vld_vec_17[16] = dep_chan_vld_16_17;
    assign in_chan_dep_data_vec_17[594 : 560] = dep_chan_data_16_17;
    assign token_in_vec_17[16] = token_16_17;
    assign in_chan_dep_vld_vec_17[17] = dep_chan_vld_18_17;
    assign in_chan_dep_data_vec_17[629 : 595] = dep_chan_data_18_17;
    assign token_in_vec_17[17] = token_18_17;
    assign in_chan_dep_vld_vec_17[18] = dep_chan_vld_33_17;
    assign in_chan_dep_data_vec_17[664 : 630] = dep_chan_data_33_17;
    assign token_in_vec_17[18] = token_33_17;
    assign dep_chan_vld_17_0 = out_chan_dep_vld_vec_17[0];
    assign dep_chan_data_17_0 = out_chan_dep_data_17;
    assign token_17_0 = token_out_vec_17[0];
    assign dep_chan_vld_17_2 = out_chan_dep_vld_vec_17[1];
    assign dep_chan_data_17_2 = out_chan_dep_data_17;
    assign token_17_2 = token_out_vec_17[1];
    assign dep_chan_vld_17_33 = out_chan_dep_vld_vec_17[2];
    assign dep_chan_data_17_33 = out_chan_dep_data_17;
    assign token_17_33 = token_out_vec_17[2];
    assign dep_chan_vld_17_1 = out_chan_dep_vld_vec_17[3];
    assign dep_chan_data_17_1 = out_chan_dep_data_17;
    assign token_17_1 = token_out_vec_17[3];
    assign dep_chan_vld_17_3 = out_chan_dep_vld_vec_17[4];
    assign dep_chan_data_17_3 = out_chan_dep_data_17;
    assign token_17_3 = token_out_vec_17[4];
    assign dep_chan_vld_17_4 = out_chan_dep_vld_vec_17[5];
    assign dep_chan_data_17_4 = out_chan_dep_data_17;
    assign token_17_4 = token_out_vec_17[5];
    assign dep_chan_vld_17_5 = out_chan_dep_vld_vec_17[6];
    assign dep_chan_data_17_5 = out_chan_dep_data_17;
    assign token_17_5 = token_out_vec_17[6];
    assign dep_chan_vld_17_6 = out_chan_dep_vld_vec_17[7];
    assign dep_chan_data_17_6 = out_chan_dep_data_17;
    assign token_17_6 = token_out_vec_17[7];
    assign dep_chan_vld_17_7 = out_chan_dep_vld_vec_17[8];
    assign dep_chan_data_17_7 = out_chan_dep_data_17;
    assign token_17_7 = token_out_vec_17[8];
    assign dep_chan_vld_17_8 = out_chan_dep_vld_vec_17[9];
    assign dep_chan_data_17_8 = out_chan_dep_data_17;
    assign token_17_8 = token_out_vec_17[9];
    assign dep_chan_vld_17_9 = out_chan_dep_vld_vec_17[10];
    assign dep_chan_data_17_9 = out_chan_dep_data_17;
    assign token_17_9 = token_out_vec_17[10];
    assign dep_chan_vld_17_10 = out_chan_dep_vld_vec_17[11];
    assign dep_chan_data_17_10 = out_chan_dep_data_17;
    assign token_17_10 = token_out_vec_17[11];
    assign dep_chan_vld_17_11 = out_chan_dep_vld_vec_17[12];
    assign dep_chan_data_17_11 = out_chan_dep_data_17;
    assign token_17_11 = token_out_vec_17[12];
    assign dep_chan_vld_17_12 = out_chan_dep_vld_vec_17[13];
    assign dep_chan_data_17_12 = out_chan_dep_data_17;
    assign token_17_12 = token_out_vec_17[13];
    assign dep_chan_vld_17_13 = out_chan_dep_vld_vec_17[14];
    assign dep_chan_data_17_13 = out_chan_dep_data_17;
    assign token_17_13 = token_out_vec_17[14];
    assign dep_chan_vld_17_14 = out_chan_dep_vld_vec_17[15];
    assign dep_chan_data_17_14 = out_chan_dep_data_17;
    assign token_17_14 = token_out_vec_17[15];
    assign dep_chan_vld_17_15 = out_chan_dep_vld_vec_17[16];
    assign dep_chan_data_17_15 = out_chan_dep_data_17;
    assign token_17_15 = token_out_vec_17[16];
    assign dep_chan_vld_17_16 = out_chan_dep_vld_vec_17[17];
    assign dep_chan_data_17_16 = out_chan_dep_data_17;
    assign token_17_16 = token_out_vec_17[17];
    assign dep_chan_vld_17_18 = out_chan_dep_vld_vec_17[18];
    assign dep_chan_data_17_18 = out_chan_dep_data_17;
    assign token_17_18 = token_out_vec_17[18];

    // Process: load_value47_U0
    kernel_pr_hls_deadlock_detect_unit #(35, 18, 19, 19) kernel_pr_hls_deadlock_detect_unit_18 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_18),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_18),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_18),
        .token_in_vec(token_in_vec_18),
        .dl_detect_in(dl_detect_out),
        .origin(origin[18]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_18),
        .out_chan_dep_data(out_chan_dep_data_18),
        .token_out_vec(token_out_vec_18),
        .dl_detect_out(dl_in_vec[18]));

    assign proc_18_data_FIFO_blk[0] = 1'b0 | (~load_value47_U0.value_r_blk_n);
    assign proc_18_data_PIPO_blk[0] = 1'b0;
    assign proc_18_start_FIFO_blk[0] = 1'b0;
    assign proc_18_TLF_FIFO_blk[0] = 1'b0;
    assign proc_18_input_sync_blk[0] = 1'b0 | (ap_sync_load_value47_U0_ap_ready & load_value47_U0.ap_idle & ~ap_sync_kernel_pr_entry98_U0_ap_ready);
    assign proc_18_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_18[0] = dl_detect_out ? proc_dep_vld_vec_18_reg[0] : (proc_18_data_FIFO_blk[0] | proc_18_data_PIPO_blk[0] | proc_18_start_FIFO_blk[0] | proc_18_TLF_FIFO_blk[0] | proc_18_input_sync_blk[0] | proc_18_output_sync_blk[0]);
    assign proc_18_data_FIFO_blk[1] = 1'b0 | (~load_value47_U0.bipedge_size_blk_n) | (~load_value47_U0.bipedge_stream_V_V15_blk_n);
    assign proc_18_data_PIPO_blk[1] = 1'b0;
    assign proc_18_start_FIFO_blk[1] = 1'b0;
    assign proc_18_TLF_FIFO_blk[1] = 1'b0;
    assign proc_18_input_sync_blk[1] = 1'b0 | (ap_sync_load_value47_U0_ap_ready & load_value47_U0.ap_idle & ~ap_sync_load_bipedge31_U0_ap_ready);
    assign proc_18_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_18[1] = dl_detect_out ? proc_dep_vld_vec_18_reg[1] : (proc_18_data_FIFO_blk[1] | proc_18_data_PIPO_blk[1] | proc_18_start_FIFO_blk[1] | proc_18_TLF_FIFO_blk[1] | proc_18_input_sync_blk[1] | proc_18_output_sync_blk[1]);
    assign proc_18_data_FIFO_blk[2] = 1'b0 | (~load_value47_U0.value_stream_V_V30_blk_n);
    assign proc_18_data_PIPO_blk[2] = 1'b0;
    assign proc_18_start_FIFO_blk[2] = 1'b0;
    assign proc_18_TLF_FIFO_blk[2] = 1'b0;
    assign proc_18_input_sync_blk[2] = 1'b0;
    assign proc_18_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_18[2] = dl_detect_out ? proc_dep_vld_vec_18_reg[2] : (proc_18_data_FIFO_blk[2] | proc_18_data_PIPO_blk[2] | proc_18_start_FIFO_blk[2] | proc_18_TLF_FIFO_blk[2] | proc_18_input_sync_blk[2] | proc_18_output_sync_blk[2]);
    assign proc_18_data_FIFO_blk[3] = 1'b0;
    assign proc_18_data_PIPO_blk[3] = 1'b0;
    assign proc_18_start_FIFO_blk[3] = 1'b0;
    assign proc_18_TLF_FIFO_blk[3] = 1'b0;
    assign proc_18_input_sync_blk[3] = 1'b0 | (ap_sync_load_value47_U0_ap_ready & load_value47_U0.ap_idle & ~ap_sync_load_bipedge30_U0_ap_ready);
    assign proc_18_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_18[3] = dl_detect_out ? proc_dep_vld_vec_18_reg[3] : (proc_18_data_FIFO_blk[3] | proc_18_data_PIPO_blk[3] | proc_18_start_FIFO_blk[3] | proc_18_TLF_FIFO_blk[3] | proc_18_input_sync_blk[3] | proc_18_output_sync_blk[3]);
    assign proc_18_data_FIFO_blk[4] = 1'b0;
    assign proc_18_data_PIPO_blk[4] = 1'b0;
    assign proc_18_start_FIFO_blk[4] = 1'b0;
    assign proc_18_TLF_FIFO_blk[4] = 1'b0;
    assign proc_18_input_sync_blk[4] = 1'b0 | (ap_sync_load_value47_U0_ap_ready & load_value47_U0.ap_idle & ~ap_sync_load_value32_U0_ap_ready);
    assign proc_18_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_18[4] = dl_detect_out ? proc_dep_vld_vec_18_reg[4] : (proc_18_data_FIFO_blk[4] | proc_18_data_PIPO_blk[4] | proc_18_start_FIFO_blk[4] | proc_18_TLF_FIFO_blk[4] | proc_18_input_sync_blk[4] | proc_18_output_sync_blk[4]);
    assign proc_18_data_FIFO_blk[5] = 1'b0;
    assign proc_18_data_PIPO_blk[5] = 1'b0;
    assign proc_18_start_FIFO_blk[5] = 1'b0;
    assign proc_18_TLF_FIFO_blk[5] = 1'b0;
    assign proc_18_input_sync_blk[5] = 1'b0 | (ap_sync_load_value47_U0_ap_ready & load_value47_U0.ap_idle & ~ap_sync_load_value33_U0_ap_ready);
    assign proc_18_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_18[5] = dl_detect_out ? proc_dep_vld_vec_18_reg[5] : (proc_18_data_FIFO_blk[5] | proc_18_data_PIPO_blk[5] | proc_18_start_FIFO_blk[5] | proc_18_TLF_FIFO_blk[5] | proc_18_input_sync_blk[5] | proc_18_output_sync_blk[5]);
    assign proc_18_data_FIFO_blk[6] = 1'b0;
    assign proc_18_data_PIPO_blk[6] = 1'b0;
    assign proc_18_start_FIFO_blk[6] = 1'b0;
    assign proc_18_TLF_FIFO_blk[6] = 1'b0;
    assign proc_18_input_sync_blk[6] = 1'b0 | (ap_sync_load_value47_U0_ap_ready & load_value47_U0.ap_idle & ~ap_sync_load_value34_U0_ap_ready);
    assign proc_18_output_sync_blk[6] = 1'b0;
    assign proc_dep_vld_vec_18[6] = dl_detect_out ? proc_dep_vld_vec_18_reg[6] : (proc_18_data_FIFO_blk[6] | proc_18_data_PIPO_blk[6] | proc_18_start_FIFO_blk[6] | proc_18_TLF_FIFO_blk[6] | proc_18_input_sync_blk[6] | proc_18_output_sync_blk[6]);
    assign proc_18_data_FIFO_blk[7] = 1'b0;
    assign proc_18_data_PIPO_blk[7] = 1'b0;
    assign proc_18_start_FIFO_blk[7] = 1'b0;
    assign proc_18_TLF_FIFO_blk[7] = 1'b0;
    assign proc_18_input_sync_blk[7] = 1'b0 | (ap_sync_load_value47_U0_ap_ready & load_value47_U0.ap_idle & ~ap_sync_load_value35_U0_ap_ready);
    assign proc_18_output_sync_blk[7] = 1'b0;
    assign proc_dep_vld_vec_18[7] = dl_detect_out ? proc_dep_vld_vec_18_reg[7] : (proc_18_data_FIFO_blk[7] | proc_18_data_PIPO_blk[7] | proc_18_start_FIFO_blk[7] | proc_18_TLF_FIFO_blk[7] | proc_18_input_sync_blk[7] | proc_18_output_sync_blk[7]);
    assign proc_18_data_FIFO_blk[8] = 1'b0;
    assign proc_18_data_PIPO_blk[8] = 1'b0;
    assign proc_18_start_FIFO_blk[8] = 1'b0;
    assign proc_18_TLF_FIFO_blk[8] = 1'b0;
    assign proc_18_input_sync_blk[8] = 1'b0 | (ap_sync_load_value47_U0_ap_ready & load_value47_U0.ap_idle & ~ap_sync_load_value36_U0_ap_ready);
    assign proc_18_output_sync_blk[8] = 1'b0;
    assign proc_dep_vld_vec_18[8] = dl_detect_out ? proc_dep_vld_vec_18_reg[8] : (proc_18_data_FIFO_blk[8] | proc_18_data_PIPO_blk[8] | proc_18_start_FIFO_blk[8] | proc_18_TLF_FIFO_blk[8] | proc_18_input_sync_blk[8] | proc_18_output_sync_blk[8]);
    assign proc_18_data_FIFO_blk[9] = 1'b0;
    assign proc_18_data_PIPO_blk[9] = 1'b0;
    assign proc_18_start_FIFO_blk[9] = 1'b0;
    assign proc_18_TLF_FIFO_blk[9] = 1'b0;
    assign proc_18_input_sync_blk[9] = 1'b0 | (ap_sync_load_value47_U0_ap_ready & load_value47_U0.ap_idle & ~ap_sync_load_value37_U0_ap_ready);
    assign proc_18_output_sync_blk[9] = 1'b0;
    assign proc_dep_vld_vec_18[9] = dl_detect_out ? proc_dep_vld_vec_18_reg[9] : (proc_18_data_FIFO_blk[9] | proc_18_data_PIPO_blk[9] | proc_18_start_FIFO_blk[9] | proc_18_TLF_FIFO_blk[9] | proc_18_input_sync_blk[9] | proc_18_output_sync_blk[9]);
    assign proc_18_data_FIFO_blk[10] = 1'b0;
    assign proc_18_data_PIPO_blk[10] = 1'b0;
    assign proc_18_start_FIFO_blk[10] = 1'b0;
    assign proc_18_TLF_FIFO_blk[10] = 1'b0;
    assign proc_18_input_sync_blk[10] = 1'b0 | (ap_sync_load_value47_U0_ap_ready & load_value47_U0.ap_idle & ~ap_sync_load_value38_U0_ap_ready);
    assign proc_18_output_sync_blk[10] = 1'b0;
    assign proc_dep_vld_vec_18[10] = dl_detect_out ? proc_dep_vld_vec_18_reg[10] : (proc_18_data_FIFO_blk[10] | proc_18_data_PIPO_blk[10] | proc_18_start_FIFO_blk[10] | proc_18_TLF_FIFO_blk[10] | proc_18_input_sync_blk[10] | proc_18_output_sync_blk[10]);
    assign proc_18_data_FIFO_blk[11] = 1'b0;
    assign proc_18_data_PIPO_blk[11] = 1'b0;
    assign proc_18_start_FIFO_blk[11] = 1'b0;
    assign proc_18_TLF_FIFO_blk[11] = 1'b0;
    assign proc_18_input_sync_blk[11] = 1'b0 | (ap_sync_load_value47_U0_ap_ready & load_value47_U0.ap_idle & ~ap_sync_load_value39_U0_ap_ready);
    assign proc_18_output_sync_blk[11] = 1'b0;
    assign proc_dep_vld_vec_18[11] = dl_detect_out ? proc_dep_vld_vec_18_reg[11] : (proc_18_data_FIFO_blk[11] | proc_18_data_PIPO_blk[11] | proc_18_start_FIFO_blk[11] | proc_18_TLF_FIFO_blk[11] | proc_18_input_sync_blk[11] | proc_18_output_sync_blk[11]);
    assign proc_18_data_FIFO_blk[12] = 1'b0;
    assign proc_18_data_PIPO_blk[12] = 1'b0;
    assign proc_18_start_FIFO_blk[12] = 1'b0;
    assign proc_18_TLF_FIFO_blk[12] = 1'b0;
    assign proc_18_input_sync_blk[12] = 1'b0 | (ap_sync_load_value47_U0_ap_ready & load_value47_U0.ap_idle & ~ap_sync_load_value40_U0_ap_ready);
    assign proc_18_output_sync_blk[12] = 1'b0;
    assign proc_dep_vld_vec_18[12] = dl_detect_out ? proc_dep_vld_vec_18_reg[12] : (proc_18_data_FIFO_blk[12] | proc_18_data_PIPO_blk[12] | proc_18_start_FIFO_blk[12] | proc_18_TLF_FIFO_blk[12] | proc_18_input_sync_blk[12] | proc_18_output_sync_blk[12]);
    assign proc_18_data_FIFO_blk[13] = 1'b0;
    assign proc_18_data_PIPO_blk[13] = 1'b0;
    assign proc_18_start_FIFO_blk[13] = 1'b0;
    assign proc_18_TLF_FIFO_blk[13] = 1'b0;
    assign proc_18_input_sync_blk[13] = 1'b0 | (ap_sync_load_value47_U0_ap_ready & load_value47_U0.ap_idle & ~ap_sync_load_value41_U0_ap_ready);
    assign proc_18_output_sync_blk[13] = 1'b0;
    assign proc_dep_vld_vec_18[13] = dl_detect_out ? proc_dep_vld_vec_18_reg[13] : (proc_18_data_FIFO_blk[13] | proc_18_data_PIPO_blk[13] | proc_18_start_FIFO_blk[13] | proc_18_TLF_FIFO_blk[13] | proc_18_input_sync_blk[13] | proc_18_output_sync_blk[13]);
    assign proc_18_data_FIFO_blk[14] = 1'b0;
    assign proc_18_data_PIPO_blk[14] = 1'b0;
    assign proc_18_start_FIFO_blk[14] = 1'b0;
    assign proc_18_TLF_FIFO_blk[14] = 1'b0;
    assign proc_18_input_sync_blk[14] = 1'b0 | (ap_sync_load_value47_U0_ap_ready & load_value47_U0.ap_idle & ~ap_sync_load_value42_U0_ap_ready);
    assign proc_18_output_sync_blk[14] = 1'b0;
    assign proc_dep_vld_vec_18[14] = dl_detect_out ? proc_dep_vld_vec_18_reg[14] : (proc_18_data_FIFO_blk[14] | proc_18_data_PIPO_blk[14] | proc_18_start_FIFO_blk[14] | proc_18_TLF_FIFO_blk[14] | proc_18_input_sync_blk[14] | proc_18_output_sync_blk[14]);
    assign proc_18_data_FIFO_blk[15] = 1'b0;
    assign proc_18_data_PIPO_blk[15] = 1'b0;
    assign proc_18_start_FIFO_blk[15] = 1'b0;
    assign proc_18_TLF_FIFO_blk[15] = 1'b0;
    assign proc_18_input_sync_blk[15] = 1'b0 | (ap_sync_load_value47_U0_ap_ready & load_value47_U0.ap_idle & ~ap_sync_load_value43_U0_ap_ready);
    assign proc_18_output_sync_blk[15] = 1'b0;
    assign proc_dep_vld_vec_18[15] = dl_detect_out ? proc_dep_vld_vec_18_reg[15] : (proc_18_data_FIFO_blk[15] | proc_18_data_PIPO_blk[15] | proc_18_start_FIFO_blk[15] | proc_18_TLF_FIFO_blk[15] | proc_18_input_sync_blk[15] | proc_18_output_sync_blk[15]);
    assign proc_18_data_FIFO_blk[16] = 1'b0;
    assign proc_18_data_PIPO_blk[16] = 1'b0;
    assign proc_18_start_FIFO_blk[16] = 1'b0;
    assign proc_18_TLF_FIFO_blk[16] = 1'b0;
    assign proc_18_input_sync_blk[16] = 1'b0 | (ap_sync_load_value47_U0_ap_ready & load_value47_U0.ap_idle & ~ap_sync_load_value44_U0_ap_ready);
    assign proc_18_output_sync_blk[16] = 1'b0;
    assign proc_dep_vld_vec_18[16] = dl_detect_out ? proc_dep_vld_vec_18_reg[16] : (proc_18_data_FIFO_blk[16] | proc_18_data_PIPO_blk[16] | proc_18_start_FIFO_blk[16] | proc_18_TLF_FIFO_blk[16] | proc_18_input_sync_blk[16] | proc_18_output_sync_blk[16]);
    assign proc_18_data_FIFO_blk[17] = 1'b0;
    assign proc_18_data_PIPO_blk[17] = 1'b0;
    assign proc_18_start_FIFO_blk[17] = 1'b0;
    assign proc_18_TLF_FIFO_blk[17] = 1'b0;
    assign proc_18_input_sync_blk[17] = 1'b0 | (ap_sync_load_value47_U0_ap_ready & load_value47_U0.ap_idle & ~ap_sync_load_value45_U0_ap_ready);
    assign proc_18_output_sync_blk[17] = 1'b0;
    assign proc_dep_vld_vec_18[17] = dl_detect_out ? proc_dep_vld_vec_18_reg[17] : (proc_18_data_FIFO_blk[17] | proc_18_data_PIPO_blk[17] | proc_18_start_FIFO_blk[17] | proc_18_TLF_FIFO_blk[17] | proc_18_input_sync_blk[17] | proc_18_output_sync_blk[17]);
    assign proc_18_data_FIFO_blk[18] = 1'b0;
    assign proc_18_data_PIPO_blk[18] = 1'b0;
    assign proc_18_start_FIFO_blk[18] = 1'b0;
    assign proc_18_TLF_FIFO_blk[18] = 1'b0;
    assign proc_18_input_sync_blk[18] = 1'b0 | (ap_sync_load_value47_U0_ap_ready & load_value47_U0.ap_idle & ~ap_sync_load_value46_U0_ap_ready);
    assign proc_18_output_sync_blk[18] = 1'b0;
    assign proc_dep_vld_vec_18[18] = dl_detect_out ? proc_dep_vld_vec_18_reg[18] : (proc_18_data_FIFO_blk[18] | proc_18_data_PIPO_blk[18] | proc_18_start_FIFO_blk[18] | proc_18_TLF_FIFO_blk[18] | proc_18_input_sync_blk[18] | proc_18_output_sync_blk[18]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_18_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_18_reg <= proc_dep_vld_vec_18;
        end
    end
    assign in_chan_dep_vld_vec_18[0] = dep_chan_vld_0_18;
    assign in_chan_dep_data_vec_18[34 : 0] = dep_chan_data_0_18;
    assign token_in_vec_18[0] = token_0_18;
    assign in_chan_dep_vld_vec_18[1] = dep_chan_vld_1_18;
    assign in_chan_dep_data_vec_18[69 : 35] = dep_chan_data_1_18;
    assign token_in_vec_18[1] = token_1_18;
    assign in_chan_dep_vld_vec_18[2] = dep_chan_vld_2_18;
    assign in_chan_dep_data_vec_18[104 : 70] = dep_chan_data_2_18;
    assign token_in_vec_18[2] = token_2_18;
    assign in_chan_dep_vld_vec_18[3] = dep_chan_vld_3_18;
    assign in_chan_dep_data_vec_18[139 : 105] = dep_chan_data_3_18;
    assign token_in_vec_18[3] = token_3_18;
    assign in_chan_dep_vld_vec_18[4] = dep_chan_vld_4_18;
    assign in_chan_dep_data_vec_18[174 : 140] = dep_chan_data_4_18;
    assign token_in_vec_18[4] = token_4_18;
    assign in_chan_dep_vld_vec_18[5] = dep_chan_vld_5_18;
    assign in_chan_dep_data_vec_18[209 : 175] = dep_chan_data_5_18;
    assign token_in_vec_18[5] = token_5_18;
    assign in_chan_dep_vld_vec_18[6] = dep_chan_vld_6_18;
    assign in_chan_dep_data_vec_18[244 : 210] = dep_chan_data_6_18;
    assign token_in_vec_18[6] = token_6_18;
    assign in_chan_dep_vld_vec_18[7] = dep_chan_vld_7_18;
    assign in_chan_dep_data_vec_18[279 : 245] = dep_chan_data_7_18;
    assign token_in_vec_18[7] = token_7_18;
    assign in_chan_dep_vld_vec_18[8] = dep_chan_vld_8_18;
    assign in_chan_dep_data_vec_18[314 : 280] = dep_chan_data_8_18;
    assign token_in_vec_18[8] = token_8_18;
    assign in_chan_dep_vld_vec_18[9] = dep_chan_vld_9_18;
    assign in_chan_dep_data_vec_18[349 : 315] = dep_chan_data_9_18;
    assign token_in_vec_18[9] = token_9_18;
    assign in_chan_dep_vld_vec_18[10] = dep_chan_vld_10_18;
    assign in_chan_dep_data_vec_18[384 : 350] = dep_chan_data_10_18;
    assign token_in_vec_18[10] = token_10_18;
    assign in_chan_dep_vld_vec_18[11] = dep_chan_vld_11_18;
    assign in_chan_dep_data_vec_18[419 : 385] = dep_chan_data_11_18;
    assign token_in_vec_18[11] = token_11_18;
    assign in_chan_dep_vld_vec_18[12] = dep_chan_vld_12_18;
    assign in_chan_dep_data_vec_18[454 : 420] = dep_chan_data_12_18;
    assign token_in_vec_18[12] = token_12_18;
    assign in_chan_dep_vld_vec_18[13] = dep_chan_vld_13_18;
    assign in_chan_dep_data_vec_18[489 : 455] = dep_chan_data_13_18;
    assign token_in_vec_18[13] = token_13_18;
    assign in_chan_dep_vld_vec_18[14] = dep_chan_vld_14_18;
    assign in_chan_dep_data_vec_18[524 : 490] = dep_chan_data_14_18;
    assign token_in_vec_18[14] = token_14_18;
    assign in_chan_dep_vld_vec_18[15] = dep_chan_vld_15_18;
    assign in_chan_dep_data_vec_18[559 : 525] = dep_chan_data_15_18;
    assign token_in_vec_18[15] = token_15_18;
    assign in_chan_dep_vld_vec_18[16] = dep_chan_vld_16_18;
    assign in_chan_dep_data_vec_18[594 : 560] = dep_chan_data_16_18;
    assign token_in_vec_18[16] = token_16_18;
    assign in_chan_dep_vld_vec_18[17] = dep_chan_vld_17_18;
    assign in_chan_dep_data_vec_18[629 : 595] = dep_chan_data_17_18;
    assign token_in_vec_18[17] = token_17_18;
    assign in_chan_dep_vld_vec_18[18] = dep_chan_vld_34_18;
    assign in_chan_dep_data_vec_18[664 : 630] = dep_chan_data_34_18;
    assign token_in_vec_18[18] = token_34_18;
    assign dep_chan_vld_18_0 = out_chan_dep_vld_vec_18[0];
    assign dep_chan_data_18_0 = out_chan_dep_data_18;
    assign token_18_0 = token_out_vec_18[0];
    assign dep_chan_vld_18_2 = out_chan_dep_vld_vec_18[1];
    assign dep_chan_data_18_2 = out_chan_dep_data_18;
    assign token_18_2 = token_out_vec_18[1];
    assign dep_chan_vld_18_34 = out_chan_dep_vld_vec_18[2];
    assign dep_chan_data_18_34 = out_chan_dep_data_18;
    assign token_18_34 = token_out_vec_18[2];
    assign dep_chan_vld_18_1 = out_chan_dep_vld_vec_18[3];
    assign dep_chan_data_18_1 = out_chan_dep_data_18;
    assign token_18_1 = token_out_vec_18[3];
    assign dep_chan_vld_18_3 = out_chan_dep_vld_vec_18[4];
    assign dep_chan_data_18_3 = out_chan_dep_data_18;
    assign token_18_3 = token_out_vec_18[4];
    assign dep_chan_vld_18_4 = out_chan_dep_vld_vec_18[5];
    assign dep_chan_data_18_4 = out_chan_dep_data_18;
    assign token_18_4 = token_out_vec_18[5];
    assign dep_chan_vld_18_5 = out_chan_dep_vld_vec_18[6];
    assign dep_chan_data_18_5 = out_chan_dep_data_18;
    assign token_18_5 = token_out_vec_18[6];
    assign dep_chan_vld_18_6 = out_chan_dep_vld_vec_18[7];
    assign dep_chan_data_18_6 = out_chan_dep_data_18;
    assign token_18_6 = token_out_vec_18[7];
    assign dep_chan_vld_18_7 = out_chan_dep_vld_vec_18[8];
    assign dep_chan_data_18_7 = out_chan_dep_data_18;
    assign token_18_7 = token_out_vec_18[8];
    assign dep_chan_vld_18_8 = out_chan_dep_vld_vec_18[9];
    assign dep_chan_data_18_8 = out_chan_dep_data_18;
    assign token_18_8 = token_out_vec_18[9];
    assign dep_chan_vld_18_9 = out_chan_dep_vld_vec_18[10];
    assign dep_chan_data_18_9 = out_chan_dep_data_18;
    assign token_18_9 = token_out_vec_18[10];
    assign dep_chan_vld_18_10 = out_chan_dep_vld_vec_18[11];
    assign dep_chan_data_18_10 = out_chan_dep_data_18;
    assign token_18_10 = token_out_vec_18[11];
    assign dep_chan_vld_18_11 = out_chan_dep_vld_vec_18[12];
    assign dep_chan_data_18_11 = out_chan_dep_data_18;
    assign token_18_11 = token_out_vec_18[12];
    assign dep_chan_vld_18_12 = out_chan_dep_vld_vec_18[13];
    assign dep_chan_data_18_12 = out_chan_dep_data_18;
    assign token_18_12 = token_out_vec_18[13];
    assign dep_chan_vld_18_13 = out_chan_dep_vld_vec_18[14];
    assign dep_chan_data_18_13 = out_chan_dep_data_18;
    assign token_18_13 = token_out_vec_18[14];
    assign dep_chan_vld_18_14 = out_chan_dep_vld_vec_18[15];
    assign dep_chan_data_18_14 = out_chan_dep_data_18;
    assign token_18_14 = token_out_vec_18[15];
    assign dep_chan_vld_18_15 = out_chan_dep_vld_vec_18[16];
    assign dep_chan_data_18_15 = out_chan_dep_data_18;
    assign token_18_15 = token_out_vec_18[16];
    assign dep_chan_vld_18_16 = out_chan_dep_vld_vec_18[17];
    assign dep_chan_data_18_16 = out_chan_dep_data_18;
    assign token_18_16 = token_out_vec_18[17];
    assign dep_chan_vld_18_17 = out_chan_dep_vld_vec_18[18];
    assign dep_chan_data_18_17 = out_chan_dep_data_18;
    assign token_18_17 = token_out_vec_18[18];

    // Process: write_back48_U0
    kernel_pr_hls_deadlock_detect_unit #(35, 19, 17, 17) kernel_pr_hls_deadlock_detect_unit_19 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_19),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_19),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_19),
        .token_in_vec(token_in_vec_19),
        .dl_detect_in(dl_detect_out),
        .origin(origin[19]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_19),
        .out_chan_dep_data(out_chan_dep_data_19),
        .token_out_vec(token_out_vec_19),
        .dl_detect_out(dl_in_vec[19]));

    assign proc_19_data_FIFO_blk[0] = 1'b0 | (~write_back48_U0.H_blk_n) | (~write_back48_U0.hyperedge_size_blk_n);
    assign proc_19_data_PIPO_blk[0] = 1'b0;
    assign proc_19_start_FIFO_blk[0] = 1'b0 | (~start_for_write_back48_U0_U.if_empty_n & write_back48_U0.ap_idle & ~start_for_write_back48_U0_U.if_write);
    assign proc_19_TLF_FIFO_blk[0] = 1'b0;
    assign proc_19_input_sync_blk[0] = 1'b0;
    assign proc_19_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_19[0] = dl_detect_out ? proc_dep_vld_vec_19_reg[0] : (proc_19_data_FIFO_blk[0] | proc_19_data_PIPO_blk[0] | proc_19_start_FIFO_blk[0] | proc_19_TLF_FIFO_blk[0] | proc_19_input_sync_blk[0] | proc_19_output_sync_blk[0]);
    assign proc_19_data_FIFO_blk[1] = 1'b0 | (~write_back48_U0.value_stream_V_V_blk_n);
    assign proc_19_data_PIPO_blk[1] = 1'b0;
    assign proc_19_start_FIFO_blk[1] = 1'b0;
    assign proc_19_TLF_FIFO_blk[1] = 1'b0;
    assign proc_19_input_sync_blk[1] = 1'b0;
    assign proc_19_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_19[1] = dl_detect_out ? proc_dep_vld_vec_19_reg[1] : (proc_19_data_FIFO_blk[1] | proc_19_data_PIPO_blk[1] | proc_19_start_FIFO_blk[1] | proc_19_TLF_FIFO_blk[1] | proc_19_input_sync_blk[1] | proc_19_output_sync_blk[1]);
    assign proc_19_data_FIFO_blk[2] = 1'b0;
    assign proc_19_data_PIPO_blk[2] = 1'b0;
    assign proc_19_start_FIFO_blk[2] = 1'b0;
    assign proc_19_TLF_FIFO_blk[2] = 1'b0;
    assign proc_19_input_sync_blk[2] = 1'b0;
    assign proc_19_output_sync_blk[2] = 1'b0 | (ap_done_reg_0 & write_back48_U0.ap_done & ~write_back49_U0.ap_done);
    assign proc_dep_vld_vec_19[2] = dl_detect_out ? proc_dep_vld_vec_19_reg[2] : (proc_19_data_FIFO_blk[2] | proc_19_data_PIPO_blk[2] | proc_19_start_FIFO_blk[2] | proc_19_TLF_FIFO_blk[2] | proc_19_input_sync_blk[2] | proc_19_output_sync_blk[2]);
    assign proc_19_data_FIFO_blk[3] = 1'b0;
    assign proc_19_data_PIPO_blk[3] = 1'b0;
    assign proc_19_start_FIFO_blk[3] = 1'b0;
    assign proc_19_TLF_FIFO_blk[3] = 1'b0;
    assign proc_19_input_sync_blk[3] = 1'b0;
    assign proc_19_output_sync_blk[3] = 1'b0 | (ap_done_reg_0 & write_back48_U0.ap_done & ~write_back50_U0.ap_done);
    assign proc_dep_vld_vec_19[3] = dl_detect_out ? proc_dep_vld_vec_19_reg[3] : (proc_19_data_FIFO_blk[3] | proc_19_data_PIPO_blk[3] | proc_19_start_FIFO_blk[3] | proc_19_TLF_FIFO_blk[3] | proc_19_input_sync_blk[3] | proc_19_output_sync_blk[3]);
    assign proc_19_data_FIFO_blk[4] = 1'b0;
    assign proc_19_data_PIPO_blk[4] = 1'b0;
    assign proc_19_start_FIFO_blk[4] = 1'b0;
    assign proc_19_TLF_FIFO_blk[4] = 1'b0;
    assign proc_19_input_sync_blk[4] = 1'b0;
    assign proc_19_output_sync_blk[4] = 1'b0 | (ap_done_reg_0 & write_back48_U0.ap_done & ~write_back51_U0.ap_done);
    assign proc_dep_vld_vec_19[4] = dl_detect_out ? proc_dep_vld_vec_19_reg[4] : (proc_19_data_FIFO_blk[4] | proc_19_data_PIPO_blk[4] | proc_19_start_FIFO_blk[4] | proc_19_TLF_FIFO_blk[4] | proc_19_input_sync_blk[4] | proc_19_output_sync_blk[4]);
    assign proc_19_data_FIFO_blk[5] = 1'b0;
    assign proc_19_data_PIPO_blk[5] = 1'b0;
    assign proc_19_start_FIFO_blk[5] = 1'b0;
    assign proc_19_TLF_FIFO_blk[5] = 1'b0;
    assign proc_19_input_sync_blk[5] = 1'b0;
    assign proc_19_output_sync_blk[5] = 1'b0 | (ap_done_reg_0 & write_back48_U0.ap_done & ~write_back52_U0.ap_done);
    assign proc_dep_vld_vec_19[5] = dl_detect_out ? proc_dep_vld_vec_19_reg[5] : (proc_19_data_FIFO_blk[5] | proc_19_data_PIPO_blk[5] | proc_19_start_FIFO_blk[5] | proc_19_TLF_FIFO_blk[5] | proc_19_input_sync_blk[5] | proc_19_output_sync_blk[5]);
    assign proc_19_data_FIFO_blk[6] = 1'b0;
    assign proc_19_data_PIPO_blk[6] = 1'b0;
    assign proc_19_start_FIFO_blk[6] = 1'b0;
    assign proc_19_TLF_FIFO_blk[6] = 1'b0;
    assign proc_19_input_sync_blk[6] = 1'b0;
    assign proc_19_output_sync_blk[6] = 1'b0 | (ap_done_reg_0 & write_back48_U0.ap_done & ~write_back53_U0.ap_done);
    assign proc_dep_vld_vec_19[6] = dl_detect_out ? proc_dep_vld_vec_19_reg[6] : (proc_19_data_FIFO_blk[6] | proc_19_data_PIPO_blk[6] | proc_19_start_FIFO_blk[6] | proc_19_TLF_FIFO_blk[6] | proc_19_input_sync_blk[6] | proc_19_output_sync_blk[6]);
    assign proc_19_data_FIFO_blk[7] = 1'b0;
    assign proc_19_data_PIPO_blk[7] = 1'b0;
    assign proc_19_start_FIFO_blk[7] = 1'b0;
    assign proc_19_TLF_FIFO_blk[7] = 1'b0;
    assign proc_19_input_sync_blk[7] = 1'b0;
    assign proc_19_output_sync_blk[7] = 1'b0 | (ap_done_reg_0 & write_back48_U0.ap_done & ~write_back54_U0.ap_done);
    assign proc_dep_vld_vec_19[7] = dl_detect_out ? proc_dep_vld_vec_19_reg[7] : (proc_19_data_FIFO_blk[7] | proc_19_data_PIPO_blk[7] | proc_19_start_FIFO_blk[7] | proc_19_TLF_FIFO_blk[7] | proc_19_input_sync_blk[7] | proc_19_output_sync_blk[7]);
    assign proc_19_data_FIFO_blk[8] = 1'b0;
    assign proc_19_data_PIPO_blk[8] = 1'b0;
    assign proc_19_start_FIFO_blk[8] = 1'b0;
    assign proc_19_TLF_FIFO_blk[8] = 1'b0;
    assign proc_19_input_sync_blk[8] = 1'b0;
    assign proc_19_output_sync_blk[8] = 1'b0 | (ap_done_reg_0 & write_back48_U0.ap_done & ~write_back55_U0.ap_done);
    assign proc_dep_vld_vec_19[8] = dl_detect_out ? proc_dep_vld_vec_19_reg[8] : (proc_19_data_FIFO_blk[8] | proc_19_data_PIPO_blk[8] | proc_19_start_FIFO_blk[8] | proc_19_TLF_FIFO_blk[8] | proc_19_input_sync_blk[8] | proc_19_output_sync_blk[8]);
    assign proc_19_data_FIFO_blk[9] = 1'b0;
    assign proc_19_data_PIPO_blk[9] = 1'b0;
    assign proc_19_start_FIFO_blk[9] = 1'b0;
    assign proc_19_TLF_FIFO_blk[9] = 1'b0;
    assign proc_19_input_sync_blk[9] = 1'b0;
    assign proc_19_output_sync_blk[9] = 1'b0 | (ap_done_reg_0 & write_back48_U0.ap_done & ~write_back56_U0.ap_done);
    assign proc_dep_vld_vec_19[9] = dl_detect_out ? proc_dep_vld_vec_19_reg[9] : (proc_19_data_FIFO_blk[9] | proc_19_data_PIPO_blk[9] | proc_19_start_FIFO_blk[9] | proc_19_TLF_FIFO_blk[9] | proc_19_input_sync_blk[9] | proc_19_output_sync_blk[9]);
    assign proc_19_data_FIFO_blk[10] = 1'b0;
    assign proc_19_data_PIPO_blk[10] = 1'b0;
    assign proc_19_start_FIFO_blk[10] = 1'b0;
    assign proc_19_TLF_FIFO_blk[10] = 1'b0;
    assign proc_19_input_sync_blk[10] = 1'b0;
    assign proc_19_output_sync_blk[10] = 1'b0 | (ap_done_reg_0 & write_back48_U0.ap_done & ~write_back57_U0.ap_done);
    assign proc_dep_vld_vec_19[10] = dl_detect_out ? proc_dep_vld_vec_19_reg[10] : (proc_19_data_FIFO_blk[10] | proc_19_data_PIPO_blk[10] | proc_19_start_FIFO_blk[10] | proc_19_TLF_FIFO_blk[10] | proc_19_input_sync_blk[10] | proc_19_output_sync_blk[10]);
    assign proc_19_data_FIFO_blk[11] = 1'b0;
    assign proc_19_data_PIPO_blk[11] = 1'b0;
    assign proc_19_start_FIFO_blk[11] = 1'b0;
    assign proc_19_TLF_FIFO_blk[11] = 1'b0;
    assign proc_19_input_sync_blk[11] = 1'b0;
    assign proc_19_output_sync_blk[11] = 1'b0 | (ap_done_reg_0 & write_back48_U0.ap_done & ~write_back58_U0.ap_done);
    assign proc_dep_vld_vec_19[11] = dl_detect_out ? proc_dep_vld_vec_19_reg[11] : (proc_19_data_FIFO_blk[11] | proc_19_data_PIPO_blk[11] | proc_19_start_FIFO_blk[11] | proc_19_TLF_FIFO_blk[11] | proc_19_input_sync_blk[11] | proc_19_output_sync_blk[11]);
    assign proc_19_data_FIFO_blk[12] = 1'b0;
    assign proc_19_data_PIPO_blk[12] = 1'b0;
    assign proc_19_start_FIFO_blk[12] = 1'b0;
    assign proc_19_TLF_FIFO_blk[12] = 1'b0;
    assign proc_19_input_sync_blk[12] = 1'b0;
    assign proc_19_output_sync_blk[12] = 1'b0 | (ap_done_reg_0 & write_back48_U0.ap_done & ~write_back59_U0.ap_done);
    assign proc_dep_vld_vec_19[12] = dl_detect_out ? proc_dep_vld_vec_19_reg[12] : (proc_19_data_FIFO_blk[12] | proc_19_data_PIPO_blk[12] | proc_19_start_FIFO_blk[12] | proc_19_TLF_FIFO_blk[12] | proc_19_input_sync_blk[12] | proc_19_output_sync_blk[12]);
    assign proc_19_data_FIFO_blk[13] = 1'b0;
    assign proc_19_data_PIPO_blk[13] = 1'b0;
    assign proc_19_start_FIFO_blk[13] = 1'b0;
    assign proc_19_TLF_FIFO_blk[13] = 1'b0;
    assign proc_19_input_sync_blk[13] = 1'b0;
    assign proc_19_output_sync_blk[13] = 1'b0 | (ap_done_reg_0 & write_back48_U0.ap_done & ~write_back60_U0.ap_done);
    assign proc_dep_vld_vec_19[13] = dl_detect_out ? proc_dep_vld_vec_19_reg[13] : (proc_19_data_FIFO_blk[13] | proc_19_data_PIPO_blk[13] | proc_19_start_FIFO_blk[13] | proc_19_TLF_FIFO_blk[13] | proc_19_input_sync_blk[13] | proc_19_output_sync_blk[13]);
    assign proc_19_data_FIFO_blk[14] = 1'b0;
    assign proc_19_data_PIPO_blk[14] = 1'b0;
    assign proc_19_start_FIFO_blk[14] = 1'b0;
    assign proc_19_TLF_FIFO_blk[14] = 1'b0;
    assign proc_19_input_sync_blk[14] = 1'b0;
    assign proc_19_output_sync_blk[14] = 1'b0 | (ap_done_reg_0 & write_back48_U0.ap_done & ~write_back61_U0.ap_done);
    assign proc_dep_vld_vec_19[14] = dl_detect_out ? proc_dep_vld_vec_19_reg[14] : (proc_19_data_FIFO_blk[14] | proc_19_data_PIPO_blk[14] | proc_19_start_FIFO_blk[14] | proc_19_TLF_FIFO_blk[14] | proc_19_input_sync_blk[14] | proc_19_output_sync_blk[14]);
    assign proc_19_data_FIFO_blk[15] = 1'b0;
    assign proc_19_data_PIPO_blk[15] = 1'b0;
    assign proc_19_start_FIFO_blk[15] = 1'b0;
    assign proc_19_TLF_FIFO_blk[15] = 1'b0;
    assign proc_19_input_sync_blk[15] = 1'b0;
    assign proc_19_output_sync_blk[15] = 1'b0 | (ap_done_reg_0 & write_back48_U0.ap_done & ~write_back62_U0.ap_done);
    assign proc_dep_vld_vec_19[15] = dl_detect_out ? proc_dep_vld_vec_19_reg[15] : (proc_19_data_FIFO_blk[15] | proc_19_data_PIPO_blk[15] | proc_19_start_FIFO_blk[15] | proc_19_TLF_FIFO_blk[15] | proc_19_input_sync_blk[15] | proc_19_output_sync_blk[15]);
    assign proc_19_data_FIFO_blk[16] = 1'b0;
    assign proc_19_data_PIPO_blk[16] = 1'b0;
    assign proc_19_start_FIFO_blk[16] = 1'b0;
    assign proc_19_TLF_FIFO_blk[16] = 1'b0;
    assign proc_19_input_sync_blk[16] = 1'b0;
    assign proc_19_output_sync_blk[16] = 1'b0 | (ap_done_reg_0 & write_back48_U0.ap_done & ~write_back63_U0.ap_done);
    assign proc_dep_vld_vec_19[16] = dl_detect_out ? proc_dep_vld_vec_19_reg[16] : (proc_19_data_FIFO_blk[16] | proc_19_data_PIPO_blk[16] | proc_19_start_FIFO_blk[16] | proc_19_TLF_FIFO_blk[16] | proc_19_input_sync_blk[16] | proc_19_output_sync_blk[16]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_19_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_19_reg <= proc_dep_vld_vec_19;
        end
    end
    assign in_chan_dep_vld_vec_19[0] = dep_chan_vld_0_19;
    assign in_chan_dep_data_vec_19[34 : 0] = dep_chan_data_0_19;
    assign token_in_vec_19[0] = token_0_19;
    assign in_chan_dep_vld_vec_19[1] = dep_chan_vld_3_19;
    assign in_chan_dep_data_vec_19[69 : 35] = dep_chan_data_3_19;
    assign token_in_vec_19[1] = token_3_19;
    assign in_chan_dep_vld_vec_19[2] = dep_chan_vld_20_19;
    assign in_chan_dep_data_vec_19[104 : 70] = dep_chan_data_20_19;
    assign token_in_vec_19[2] = token_20_19;
    assign in_chan_dep_vld_vec_19[3] = dep_chan_vld_21_19;
    assign in_chan_dep_data_vec_19[139 : 105] = dep_chan_data_21_19;
    assign token_in_vec_19[3] = token_21_19;
    assign in_chan_dep_vld_vec_19[4] = dep_chan_vld_22_19;
    assign in_chan_dep_data_vec_19[174 : 140] = dep_chan_data_22_19;
    assign token_in_vec_19[4] = token_22_19;
    assign in_chan_dep_vld_vec_19[5] = dep_chan_vld_23_19;
    assign in_chan_dep_data_vec_19[209 : 175] = dep_chan_data_23_19;
    assign token_in_vec_19[5] = token_23_19;
    assign in_chan_dep_vld_vec_19[6] = dep_chan_vld_24_19;
    assign in_chan_dep_data_vec_19[244 : 210] = dep_chan_data_24_19;
    assign token_in_vec_19[6] = token_24_19;
    assign in_chan_dep_vld_vec_19[7] = dep_chan_vld_25_19;
    assign in_chan_dep_data_vec_19[279 : 245] = dep_chan_data_25_19;
    assign token_in_vec_19[7] = token_25_19;
    assign in_chan_dep_vld_vec_19[8] = dep_chan_vld_26_19;
    assign in_chan_dep_data_vec_19[314 : 280] = dep_chan_data_26_19;
    assign token_in_vec_19[8] = token_26_19;
    assign in_chan_dep_vld_vec_19[9] = dep_chan_vld_27_19;
    assign in_chan_dep_data_vec_19[349 : 315] = dep_chan_data_27_19;
    assign token_in_vec_19[9] = token_27_19;
    assign in_chan_dep_vld_vec_19[10] = dep_chan_vld_28_19;
    assign in_chan_dep_data_vec_19[384 : 350] = dep_chan_data_28_19;
    assign token_in_vec_19[10] = token_28_19;
    assign in_chan_dep_vld_vec_19[11] = dep_chan_vld_29_19;
    assign in_chan_dep_data_vec_19[419 : 385] = dep_chan_data_29_19;
    assign token_in_vec_19[11] = token_29_19;
    assign in_chan_dep_vld_vec_19[12] = dep_chan_vld_30_19;
    assign in_chan_dep_data_vec_19[454 : 420] = dep_chan_data_30_19;
    assign token_in_vec_19[12] = token_30_19;
    assign in_chan_dep_vld_vec_19[13] = dep_chan_vld_31_19;
    assign in_chan_dep_data_vec_19[489 : 455] = dep_chan_data_31_19;
    assign token_in_vec_19[13] = token_31_19;
    assign in_chan_dep_vld_vec_19[14] = dep_chan_vld_32_19;
    assign in_chan_dep_data_vec_19[524 : 490] = dep_chan_data_32_19;
    assign token_in_vec_19[14] = token_32_19;
    assign in_chan_dep_vld_vec_19[15] = dep_chan_vld_33_19;
    assign in_chan_dep_data_vec_19[559 : 525] = dep_chan_data_33_19;
    assign token_in_vec_19[15] = token_33_19;
    assign in_chan_dep_vld_vec_19[16] = dep_chan_vld_34_19;
    assign in_chan_dep_data_vec_19[594 : 560] = dep_chan_data_34_19;
    assign token_in_vec_19[16] = token_34_19;
    assign dep_chan_vld_19_0 = out_chan_dep_vld_vec_19[0];
    assign dep_chan_data_19_0 = out_chan_dep_data_19;
    assign token_19_0 = token_out_vec_19[0];
    assign dep_chan_vld_19_3 = out_chan_dep_vld_vec_19[1];
    assign dep_chan_data_19_3 = out_chan_dep_data_19;
    assign token_19_3 = token_out_vec_19[1];
    assign dep_chan_vld_19_20 = out_chan_dep_vld_vec_19[2];
    assign dep_chan_data_19_20 = out_chan_dep_data_19;
    assign token_19_20 = token_out_vec_19[2];
    assign dep_chan_vld_19_21 = out_chan_dep_vld_vec_19[3];
    assign dep_chan_data_19_21 = out_chan_dep_data_19;
    assign token_19_21 = token_out_vec_19[3];
    assign dep_chan_vld_19_22 = out_chan_dep_vld_vec_19[4];
    assign dep_chan_data_19_22 = out_chan_dep_data_19;
    assign token_19_22 = token_out_vec_19[4];
    assign dep_chan_vld_19_23 = out_chan_dep_vld_vec_19[5];
    assign dep_chan_data_19_23 = out_chan_dep_data_19;
    assign token_19_23 = token_out_vec_19[5];
    assign dep_chan_vld_19_24 = out_chan_dep_vld_vec_19[6];
    assign dep_chan_data_19_24 = out_chan_dep_data_19;
    assign token_19_24 = token_out_vec_19[6];
    assign dep_chan_vld_19_25 = out_chan_dep_vld_vec_19[7];
    assign dep_chan_data_19_25 = out_chan_dep_data_19;
    assign token_19_25 = token_out_vec_19[7];
    assign dep_chan_vld_19_26 = out_chan_dep_vld_vec_19[8];
    assign dep_chan_data_19_26 = out_chan_dep_data_19;
    assign token_19_26 = token_out_vec_19[8];
    assign dep_chan_vld_19_27 = out_chan_dep_vld_vec_19[9];
    assign dep_chan_data_19_27 = out_chan_dep_data_19;
    assign token_19_27 = token_out_vec_19[9];
    assign dep_chan_vld_19_28 = out_chan_dep_vld_vec_19[10];
    assign dep_chan_data_19_28 = out_chan_dep_data_19;
    assign token_19_28 = token_out_vec_19[10];
    assign dep_chan_vld_19_29 = out_chan_dep_vld_vec_19[11];
    assign dep_chan_data_19_29 = out_chan_dep_data_19;
    assign token_19_29 = token_out_vec_19[11];
    assign dep_chan_vld_19_30 = out_chan_dep_vld_vec_19[12];
    assign dep_chan_data_19_30 = out_chan_dep_data_19;
    assign token_19_30 = token_out_vec_19[12];
    assign dep_chan_vld_19_31 = out_chan_dep_vld_vec_19[13];
    assign dep_chan_data_19_31 = out_chan_dep_data_19;
    assign token_19_31 = token_out_vec_19[13];
    assign dep_chan_vld_19_32 = out_chan_dep_vld_vec_19[14];
    assign dep_chan_data_19_32 = out_chan_dep_data_19;
    assign token_19_32 = token_out_vec_19[14];
    assign dep_chan_vld_19_33 = out_chan_dep_vld_vec_19[15];
    assign dep_chan_data_19_33 = out_chan_dep_data_19;
    assign token_19_33 = token_out_vec_19[15];
    assign dep_chan_vld_19_34 = out_chan_dep_vld_vec_19[16];
    assign dep_chan_data_19_34 = out_chan_dep_data_19;
    assign token_19_34 = token_out_vec_19[16];

    // Process: write_back49_U0
    kernel_pr_hls_deadlock_detect_unit #(35, 20, 17, 17) kernel_pr_hls_deadlock_detect_unit_20 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_20),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_20),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_20),
        .token_in_vec(token_in_vec_20),
        .dl_detect_in(dl_detect_out),
        .origin(origin[20]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_20),
        .out_chan_dep_data(out_chan_dep_data_20),
        .token_out_vec(token_out_vec_20),
        .dl_detect_out(dl_in_vec[20]));

    assign proc_20_data_FIFO_blk[0] = 1'b0 | (~write_back49_U0.H_blk_n) | (~write_back49_U0.hyperedge_size_blk_n);
    assign proc_20_data_PIPO_blk[0] = 1'b0;
    assign proc_20_start_FIFO_blk[0] = 1'b0 | (~start_for_write_back49_U0_U.if_empty_n & write_back49_U0.ap_idle & ~start_for_write_back49_U0_U.if_write);
    assign proc_20_TLF_FIFO_blk[0] = 1'b0;
    assign proc_20_input_sync_blk[0] = 1'b0;
    assign proc_20_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_20[0] = dl_detect_out ? proc_dep_vld_vec_20_reg[0] : (proc_20_data_FIFO_blk[0] | proc_20_data_PIPO_blk[0] | proc_20_start_FIFO_blk[0] | proc_20_TLF_FIFO_blk[0] | proc_20_input_sync_blk[0] | proc_20_output_sync_blk[0]);
    assign proc_20_data_FIFO_blk[1] = 1'b0 | (~write_back49_U0.value_stream_V_V1_blk_n);
    assign proc_20_data_PIPO_blk[1] = 1'b0;
    assign proc_20_start_FIFO_blk[1] = 1'b0;
    assign proc_20_TLF_FIFO_blk[1] = 1'b0;
    assign proc_20_input_sync_blk[1] = 1'b0;
    assign proc_20_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_20[1] = dl_detect_out ? proc_dep_vld_vec_20_reg[1] : (proc_20_data_FIFO_blk[1] | proc_20_data_PIPO_blk[1] | proc_20_start_FIFO_blk[1] | proc_20_TLF_FIFO_blk[1] | proc_20_input_sync_blk[1] | proc_20_output_sync_blk[1]);
    assign proc_20_data_FIFO_blk[2] = 1'b0;
    assign proc_20_data_PIPO_blk[2] = 1'b0;
    assign proc_20_start_FIFO_blk[2] = 1'b0;
    assign proc_20_TLF_FIFO_blk[2] = 1'b0;
    assign proc_20_input_sync_blk[2] = 1'b0;
    assign proc_20_output_sync_blk[2] = 1'b0 | (ap_done_reg_1 & write_back49_U0.ap_done & ~write_back48_U0.ap_done);
    assign proc_dep_vld_vec_20[2] = dl_detect_out ? proc_dep_vld_vec_20_reg[2] : (proc_20_data_FIFO_blk[2] | proc_20_data_PIPO_blk[2] | proc_20_start_FIFO_blk[2] | proc_20_TLF_FIFO_blk[2] | proc_20_input_sync_blk[2] | proc_20_output_sync_blk[2]);
    assign proc_20_data_FIFO_blk[3] = 1'b0;
    assign proc_20_data_PIPO_blk[3] = 1'b0;
    assign proc_20_start_FIFO_blk[3] = 1'b0;
    assign proc_20_TLF_FIFO_blk[3] = 1'b0;
    assign proc_20_input_sync_blk[3] = 1'b0;
    assign proc_20_output_sync_blk[3] = 1'b0 | (ap_done_reg_1 & write_back49_U0.ap_done & ~write_back50_U0.ap_done);
    assign proc_dep_vld_vec_20[3] = dl_detect_out ? proc_dep_vld_vec_20_reg[3] : (proc_20_data_FIFO_blk[3] | proc_20_data_PIPO_blk[3] | proc_20_start_FIFO_blk[3] | proc_20_TLF_FIFO_blk[3] | proc_20_input_sync_blk[3] | proc_20_output_sync_blk[3]);
    assign proc_20_data_FIFO_blk[4] = 1'b0;
    assign proc_20_data_PIPO_blk[4] = 1'b0;
    assign proc_20_start_FIFO_blk[4] = 1'b0;
    assign proc_20_TLF_FIFO_blk[4] = 1'b0;
    assign proc_20_input_sync_blk[4] = 1'b0;
    assign proc_20_output_sync_blk[4] = 1'b0 | (ap_done_reg_1 & write_back49_U0.ap_done & ~write_back51_U0.ap_done);
    assign proc_dep_vld_vec_20[4] = dl_detect_out ? proc_dep_vld_vec_20_reg[4] : (proc_20_data_FIFO_blk[4] | proc_20_data_PIPO_blk[4] | proc_20_start_FIFO_blk[4] | proc_20_TLF_FIFO_blk[4] | proc_20_input_sync_blk[4] | proc_20_output_sync_blk[4]);
    assign proc_20_data_FIFO_blk[5] = 1'b0;
    assign proc_20_data_PIPO_blk[5] = 1'b0;
    assign proc_20_start_FIFO_blk[5] = 1'b0;
    assign proc_20_TLF_FIFO_blk[5] = 1'b0;
    assign proc_20_input_sync_blk[5] = 1'b0;
    assign proc_20_output_sync_blk[5] = 1'b0 | (ap_done_reg_1 & write_back49_U0.ap_done & ~write_back52_U0.ap_done);
    assign proc_dep_vld_vec_20[5] = dl_detect_out ? proc_dep_vld_vec_20_reg[5] : (proc_20_data_FIFO_blk[5] | proc_20_data_PIPO_blk[5] | proc_20_start_FIFO_blk[5] | proc_20_TLF_FIFO_blk[5] | proc_20_input_sync_blk[5] | proc_20_output_sync_blk[5]);
    assign proc_20_data_FIFO_blk[6] = 1'b0;
    assign proc_20_data_PIPO_blk[6] = 1'b0;
    assign proc_20_start_FIFO_blk[6] = 1'b0;
    assign proc_20_TLF_FIFO_blk[6] = 1'b0;
    assign proc_20_input_sync_blk[6] = 1'b0;
    assign proc_20_output_sync_blk[6] = 1'b0 | (ap_done_reg_1 & write_back49_U0.ap_done & ~write_back53_U0.ap_done);
    assign proc_dep_vld_vec_20[6] = dl_detect_out ? proc_dep_vld_vec_20_reg[6] : (proc_20_data_FIFO_blk[6] | proc_20_data_PIPO_blk[6] | proc_20_start_FIFO_blk[6] | proc_20_TLF_FIFO_blk[6] | proc_20_input_sync_blk[6] | proc_20_output_sync_blk[6]);
    assign proc_20_data_FIFO_blk[7] = 1'b0;
    assign proc_20_data_PIPO_blk[7] = 1'b0;
    assign proc_20_start_FIFO_blk[7] = 1'b0;
    assign proc_20_TLF_FIFO_blk[7] = 1'b0;
    assign proc_20_input_sync_blk[7] = 1'b0;
    assign proc_20_output_sync_blk[7] = 1'b0 | (ap_done_reg_1 & write_back49_U0.ap_done & ~write_back54_U0.ap_done);
    assign proc_dep_vld_vec_20[7] = dl_detect_out ? proc_dep_vld_vec_20_reg[7] : (proc_20_data_FIFO_blk[7] | proc_20_data_PIPO_blk[7] | proc_20_start_FIFO_blk[7] | proc_20_TLF_FIFO_blk[7] | proc_20_input_sync_blk[7] | proc_20_output_sync_blk[7]);
    assign proc_20_data_FIFO_blk[8] = 1'b0;
    assign proc_20_data_PIPO_blk[8] = 1'b0;
    assign proc_20_start_FIFO_blk[8] = 1'b0;
    assign proc_20_TLF_FIFO_blk[8] = 1'b0;
    assign proc_20_input_sync_blk[8] = 1'b0;
    assign proc_20_output_sync_blk[8] = 1'b0 | (ap_done_reg_1 & write_back49_U0.ap_done & ~write_back55_U0.ap_done);
    assign proc_dep_vld_vec_20[8] = dl_detect_out ? proc_dep_vld_vec_20_reg[8] : (proc_20_data_FIFO_blk[8] | proc_20_data_PIPO_blk[8] | proc_20_start_FIFO_blk[8] | proc_20_TLF_FIFO_blk[8] | proc_20_input_sync_blk[8] | proc_20_output_sync_blk[8]);
    assign proc_20_data_FIFO_blk[9] = 1'b0;
    assign proc_20_data_PIPO_blk[9] = 1'b0;
    assign proc_20_start_FIFO_blk[9] = 1'b0;
    assign proc_20_TLF_FIFO_blk[9] = 1'b0;
    assign proc_20_input_sync_blk[9] = 1'b0;
    assign proc_20_output_sync_blk[9] = 1'b0 | (ap_done_reg_1 & write_back49_U0.ap_done & ~write_back56_U0.ap_done);
    assign proc_dep_vld_vec_20[9] = dl_detect_out ? proc_dep_vld_vec_20_reg[9] : (proc_20_data_FIFO_blk[9] | proc_20_data_PIPO_blk[9] | proc_20_start_FIFO_blk[9] | proc_20_TLF_FIFO_blk[9] | proc_20_input_sync_blk[9] | proc_20_output_sync_blk[9]);
    assign proc_20_data_FIFO_blk[10] = 1'b0;
    assign proc_20_data_PIPO_blk[10] = 1'b0;
    assign proc_20_start_FIFO_blk[10] = 1'b0;
    assign proc_20_TLF_FIFO_blk[10] = 1'b0;
    assign proc_20_input_sync_blk[10] = 1'b0;
    assign proc_20_output_sync_blk[10] = 1'b0 | (ap_done_reg_1 & write_back49_U0.ap_done & ~write_back57_U0.ap_done);
    assign proc_dep_vld_vec_20[10] = dl_detect_out ? proc_dep_vld_vec_20_reg[10] : (proc_20_data_FIFO_blk[10] | proc_20_data_PIPO_blk[10] | proc_20_start_FIFO_blk[10] | proc_20_TLF_FIFO_blk[10] | proc_20_input_sync_blk[10] | proc_20_output_sync_blk[10]);
    assign proc_20_data_FIFO_blk[11] = 1'b0;
    assign proc_20_data_PIPO_blk[11] = 1'b0;
    assign proc_20_start_FIFO_blk[11] = 1'b0;
    assign proc_20_TLF_FIFO_blk[11] = 1'b0;
    assign proc_20_input_sync_blk[11] = 1'b0;
    assign proc_20_output_sync_blk[11] = 1'b0 | (ap_done_reg_1 & write_back49_U0.ap_done & ~write_back58_U0.ap_done);
    assign proc_dep_vld_vec_20[11] = dl_detect_out ? proc_dep_vld_vec_20_reg[11] : (proc_20_data_FIFO_blk[11] | proc_20_data_PIPO_blk[11] | proc_20_start_FIFO_blk[11] | proc_20_TLF_FIFO_blk[11] | proc_20_input_sync_blk[11] | proc_20_output_sync_blk[11]);
    assign proc_20_data_FIFO_blk[12] = 1'b0;
    assign proc_20_data_PIPO_blk[12] = 1'b0;
    assign proc_20_start_FIFO_blk[12] = 1'b0;
    assign proc_20_TLF_FIFO_blk[12] = 1'b0;
    assign proc_20_input_sync_blk[12] = 1'b0;
    assign proc_20_output_sync_blk[12] = 1'b0 | (ap_done_reg_1 & write_back49_U0.ap_done & ~write_back59_U0.ap_done);
    assign proc_dep_vld_vec_20[12] = dl_detect_out ? proc_dep_vld_vec_20_reg[12] : (proc_20_data_FIFO_blk[12] | proc_20_data_PIPO_blk[12] | proc_20_start_FIFO_blk[12] | proc_20_TLF_FIFO_blk[12] | proc_20_input_sync_blk[12] | proc_20_output_sync_blk[12]);
    assign proc_20_data_FIFO_blk[13] = 1'b0;
    assign proc_20_data_PIPO_blk[13] = 1'b0;
    assign proc_20_start_FIFO_blk[13] = 1'b0;
    assign proc_20_TLF_FIFO_blk[13] = 1'b0;
    assign proc_20_input_sync_blk[13] = 1'b0;
    assign proc_20_output_sync_blk[13] = 1'b0 | (ap_done_reg_1 & write_back49_U0.ap_done & ~write_back60_U0.ap_done);
    assign proc_dep_vld_vec_20[13] = dl_detect_out ? proc_dep_vld_vec_20_reg[13] : (proc_20_data_FIFO_blk[13] | proc_20_data_PIPO_blk[13] | proc_20_start_FIFO_blk[13] | proc_20_TLF_FIFO_blk[13] | proc_20_input_sync_blk[13] | proc_20_output_sync_blk[13]);
    assign proc_20_data_FIFO_blk[14] = 1'b0;
    assign proc_20_data_PIPO_blk[14] = 1'b0;
    assign proc_20_start_FIFO_blk[14] = 1'b0;
    assign proc_20_TLF_FIFO_blk[14] = 1'b0;
    assign proc_20_input_sync_blk[14] = 1'b0;
    assign proc_20_output_sync_blk[14] = 1'b0 | (ap_done_reg_1 & write_back49_U0.ap_done & ~write_back61_U0.ap_done);
    assign proc_dep_vld_vec_20[14] = dl_detect_out ? proc_dep_vld_vec_20_reg[14] : (proc_20_data_FIFO_blk[14] | proc_20_data_PIPO_blk[14] | proc_20_start_FIFO_blk[14] | proc_20_TLF_FIFO_blk[14] | proc_20_input_sync_blk[14] | proc_20_output_sync_blk[14]);
    assign proc_20_data_FIFO_blk[15] = 1'b0;
    assign proc_20_data_PIPO_blk[15] = 1'b0;
    assign proc_20_start_FIFO_blk[15] = 1'b0;
    assign proc_20_TLF_FIFO_blk[15] = 1'b0;
    assign proc_20_input_sync_blk[15] = 1'b0;
    assign proc_20_output_sync_blk[15] = 1'b0 | (ap_done_reg_1 & write_back49_U0.ap_done & ~write_back62_U0.ap_done);
    assign proc_dep_vld_vec_20[15] = dl_detect_out ? proc_dep_vld_vec_20_reg[15] : (proc_20_data_FIFO_blk[15] | proc_20_data_PIPO_blk[15] | proc_20_start_FIFO_blk[15] | proc_20_TLF_FIFO_blk[15] | proc_20_input_sync_blk[15] | proc_20_output_sync_blk[15]);
    assign proc_20_data_FIFO_blk[16] = 1'b0;
    assign proc_20_data_PIPO_blk[16] = 1'b0;
    assign proc_20_start_FIFO_blk[16] = 1'b0;
    assign proc_20_TLF_FIFO_blk[16] = 1'b0;
    assign proc_20_input_sync_blk[16] = 1'b0;
    assign proc_20_output_sync_blk[16] = 1'b0 | (ap_done_reg_1 & write_back49_U0.ap_done & ~write_back63_U0.ap_done);
    assign proc_dep_vld_vec_20[16] = dl_detect_out ? proc_dep_vld_vec_20_reg[16] : (proc_20_data_FIFO_blk[16] | proc_20_data_PIPO_blk[16] | proc_20_start_FIFO_blk[16] | proc_20_TLF_FIFO_blk[16] | proc_20_input_sync_blk[16] | proc_20_output_sync_blk[16]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_20_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_20_reg <= proc_dep_vld_vec_20;
        end
    end
    assign in_chan_dep_vld_vec_20[0] = dep_chan_vld_0_20;
    assign in_chan_dep_data_vec_20[34 : 0] = dep_chan_data_0_20;
    assign token_in_vec_20[0] = token_0_20;
    assign in_chan_dep_vld_vec_20[1] = dep_chan_vld_4_20;
    assign in_chan_dep_data_vec_20[69 : 35] = dep_chan_data_4_20;
    assign token_in_vec_20[1] = token_4_20;
    assign in_chan_dep_vld_vec_20[2] = dep_chan_vld_19_20;
    assign in_chan_dep_data_vec_20[104 : 70] = dep_chan_data_19_20;
    assign token_in_vec_20[2] = token_19_20;
    assign in_chan_dep_vld_vec_20[3] = dep_chan_vld_21_20;
    assign in_chan_dep_data_vec_20[139 : 105] = dep_chan_data_21_20;
    assign token_in_vec_20[3] = token_21_20;
    assign in_chan_dep_vld_vec_20[4] = dep_chan_vld_22_20;
    assign in_chan_dep_data_vec_20[174 : 140] = dep_chan_data_22_20;
    assign token_in_vec_20[4] = token_22_20;
    assign in_chan_dep_vld_vec_20[5] = dep_chan_vld_23_20;
    assign in_chan_dep_data_vec_20[209 : 175] = dep_chan_data_23_20;
    assign token_in_vec_20[5] = token_23_20;
    assign in_chan_dep_vld_vec_20[6] = dep_chan_vld_24_20;
    assign in_chan_dep_data_vec_20[244 : 210] = dep_chan_data_24_20;
    assign token_in_vec_20[6] = token_24_20;
    assign in_chan_dep_vld_vec_20[7] = dep_chan_vld_25_20;
    assign in_chan_dep_data_vec_20[279 : 245] = dep_chan_data_25_20;
    assign token_in_vec_20[7] = token_25_20;
    assign in_chan_dep_vld_vec_20[8] = dep_chan_vld_26_20;
    assign in_chan_dep_data_vec_20[314 : 280] = dep_chan_data_26_20;
    assign token_in_vec_20[8] = token_26_20;
    assign in_chan_dep_vld_vec_20[9] = dep_chan_vld_27_20;
    assign in_chan_dep_data_vec_20[349 : 315] = dep_chan_data_27_20;
    assign token_in_vec_20[9] = token_27_20;
    assign in_chan_dep_vld_vec_20[10] = dep_chan_vld_28_20;
    assign in_chan_dep_data_vec_20[384 : 350] = dep_chan_data_28_20;
    assign token_in_vec_20[10] = token_28_20;
    assign in_chan_dep_vld_vec_20[11] = dep_chan_vld_29_20;
    assign in_chan_dep_data_vec_20[419 : 385] = dep_chan_data_29_20;
    assign token_in_vec_20[11] = token_29_20;
    assign in_chan_dep_vld_vec_20[12] = dep_chan_vld_30_20;
    assign in_chan_dep_data_vec_20[454 : 420] = dep_chan_data_30_20;
    assign token_in_vec_20[12] = token_30_20;
    assign in_chan_dep_vld_vec_20[13] = dep_chan_vld_31_20;
    assign in_chan_dep_data_vec_20[489 : 455] = dep_chan_data_31_20;
    assign token_in_vec_20[13] = token_31_20;
    assign in_chan_dep_vld_vec_20[14] = dep_chan_vld_32_20;
    assign in_chan_dep_data_vec_20[524 : 490] = dep_chan_data_32_20;
    assign token_in_vec_20[14] = token_32_20;
    assign in_chan_dep_vld_vec_20[15] = dep_chan_vld_33_20;
    assign in_chan_dep_data_vec_20[559 : 525] = dep_chan_data_33_20;
    assign token_in_vec_20[15] = token_33_20;
    assign in_chan_dep_vld_vec_20[16] = dep_chan_vld_34_20;
    assign in_chan_dep_data_vec_20[594 : 560] = dep_chan_data_34_20;
    assign token_in_vec_20[16] = token_34_20;
    assign dep_chan_vld_20_0 = out_chan_dep_vld_vec_20[0];
    assign dep_chan_data_20_0 = out_chan_dep_data_20;
    assign token_20_0 = token_out_vec_20[0];
    assign dep_chan_vld_20_4 = out_chan_dep_vld_vec_20[1];
    assign dep_chan_data_20_4 = out_chan_dep_data_20;
    assign token_20_4 = token_out_vec_20[1];
    assign dep_chan_vld_20_19 = out_chan_dep_vld_vec_20[2];
    assign dep_chan_data_20_19 = out_chan_dep_data_20;
    assign token_20_19 = token_out_vec_20[2];
    assign dep_chan_vld_20_21 = out_chan_dep_vld_vec_20[3];
    assign dep_chan_data_20_21 = out_chan_dep_data_20;
    assign token_20_21 = token_out_vec_20[3];
    assign dep_chan_vld_20_22 = out_chan_dep_vld_vec_20[4];
    assign dep_chan_data_20_22 = out_chan_dep_data_20;
    assign token_20_22 = token_out_vec_20[4];
    assign dep_chan_vld_20_23 = out_chan_dep_vld_vec_20[5];
    assign dep_chan_data_20_23 = out_chan_dep_data_20;
    assign token_20_23 = token_out_vec_20[5];
    assign dep_chan_vld_20_24 = out_chan_dep_vld_vec_20[6];
    assign dep_chan_data_20_24 = out_chan_dep_data_20;
    assign token_20_24 = token_out_vec_20[6];
    assign dep_chan_vld_20_25 = out_chan_dep_vld_vec_20[7];
    assign dep_chan_data_20_25 = out_chan_dep_data_20;
    assign token_20_25 = token_out_vec_20[7];
    assign dep_chan_vld_20_26 = out_chan_dep_vld_vec_20[8];
    assign dep_chan_data_20_26 = out_chan_dep_data_20;
    assign token_20_26 = token_out_vec_20[8];
    assign dep_chan_vld_20_27 = out_chan_dep_vld_vec_20[9];
    assign dep_chan_data_20_27 = out_chan_dep_data_20;
    assign token_20_27 = token_out_vec_20[9];
    assign dep_chan_vld_20_28 = out_chan_dep_vld_vec_20[10];
    assign dep_chan_data_20_28 = out_chan_dep_data_20;
    assign token_20_28 = token_out_vec_20[10];
    assign dep_chan_vld_20_29 = out_chan_dep_vld_vec_20[11];
    assign dep_chan_data_20_29 = out_chan_dep_data_20;
    assign token_20_29 = token_out_vec_20[11];
    assign dep_chan_vld_20_30 = out_chan_dep_vld_vec_20[12];
    assign dep_chan_data_20_30 = out_chan_dep_data_20;
    assign token_20_30 = token_out_vec_20[12];
    assign dep_chan_vld_20_31 = out_chan_dep_vld_vec_20[13];
    assign dep_chan_data_20_31 = out_chan_dep_data_20;
    assign token_20_31 = token_out_vec_20[13];
    assign dep_chan_vld_20_32 = out_chan_dep_vld_vec_20[14];
    assign dep_chan_data_20_32 = out_chan_dep_data_20;
    assign token_20_32 = token_out_vec_20[14];
    assign dep_chan_vld_20_33 = out_chan_dep_vld_vec_20[15];
    assign dep_chan_data_20_33 = out_chan_dep_data_20;
    assign token_20_33 = token_out_vec_20[15];
    assign dep_chan_vld_20_34 = out_chan_dep_vld_vec_20[16];
    assign dep_chan_data_20_34 = out_chan_dep_data_20;
    assign token_20_34 = token_out_vec_20[16];

    // Process: write_back50_U0
    kernel_pr_hls_deadlock_detect_unit #(35, 21, 17, 17) kernel_pr_hls_deadlock_detect_unit_21 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_21),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_21),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_21),
        .token_in_vec(token_in_vec_21),
        .dl_detect_in(dl_detect_out),
        .origin(origin[21]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_21),
        .out_chan_dep_data(out_chan_dep_data_21),
        .token_out_vec(token_out_vec_21),
        .dl_detect_out(dl_in_vec[21]));

    assign proc_21_data_FIFO_blk[0] = 1'b0 | (~write_back50_U0.H_blk_n) | (~write_back50_U0.hyperedge_size_blk_n);
    assign proc_21_data_PIPO_blk[0] = 1'b0;
    assign proc_21_start_FIFO_blk[0] = 1'b0 | (~start_for_write_back50_U0_U.if_empty_n & write_back50_U0.ap_idle & ~start_for_write_back50_U0_U.if_write);
    assign proc_21_TLF_FIFO_blk[0] = 1'b0;
    assign proc_21_input_sync_blk[0] = 1'b0;
    assign proc_21_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_21[0] = dl_detect_out ? proc_dep_vld_vec_21_reg[0] : (proc_21_data_FIFO_blk[0] | proc_21_data_PIPO_blk[0] | proc_21_start_FIFO_blk[0] | proc_21_TLF_FIFO_blk[0] | proc_21_input_sync_blk[0] | proc_21_output_sync_blk[0]);
    assign proc_21_data_FIFO_blk[1] = 1'b0 | (~write_back50_U0.value_stream_V_V2_blk_n);
    assign proc_21_data_PIPO_blk[1] = 1'b0;
    assign proc_21_start_FIFO_blk[1] = 1'b0;
    assign proc_21_TLF_FIFO_blk[1] = 1'b0;
    assign proc_21_input_sync_blk[1] = 1'b0;
    assign proc_21_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_21[1] = dl_detect_out ? proc_dep_vld_vec_21_reg[1] : (proc_21_data_FIFO_blk[1] | proc_21_data_PIPO_blk[1] | proc_21_start_FIFO_blk[1] | proc_21_TLF_FIFO_blk[1] | proc_21_input_sync_blk[1] | proc_21_output_sync_blk[1]);
    assign proc_21_data_FIFO_blk[2] = 1'b0;
    assign proc_21_data_PIPO_blk[2] = 1'b0;
    assign proc_21_start_FIFO_blk[2] = 1'b0;
    assign proc_21_TLF_FIFO_blk[2] = 1'b0;
    assign proc_21_input_sync_blk[2] = 1'b0;
    assign proc_21_output_sync_blk[2] = 1'b0 | (ap_done_reg_2 & write_back50_U0.ap_done & ~write_back48_U0.ap_done);
    assign proc_dep_vld_vec_21[2] = dl_detect_out ? proc_dep_vld_vec_21_reg[2] : (proc_21_data_FIFO_blk[2] | proc_21_data_PIPO_blk[2] | proc_21_start_FIFO_blk[2] | proc_21_TLF_FIFO_blk[2] | proc_21_input_sync_blk[2] | proc_21_output_sync_blk[2]);
    assign proc_21_data_FIFO_blk[3] = 1'b0;
    assign proc_21_data_PIPO_blk[3] = 1'b0;
    assign proc_21_start_FIFO_blk[3] = 1'b0;
    assign proc_21_TLF_FIFO_blk[3] = 1'b0;
    assign proc_21_input_sync_blk[3] = 1'b0;
    assign proc_21_output_sync_blk[3] = 1'b0 | (ap_done_reg_2 & write_back50_U0.ap_done & ~write_back49_U0.ap_done);
    assign proc_dep_vld_vec_21[3] = dl_detect_out ? proc_dep_vld_vec_21_reg[3] : (proc_21_data_FIFO_blk[3] | proc_21_data_PIPO_blk[3] | proc_21_start_FIFO_blk[3] | proc_21_TLF_FIFO_blk[3] | proc_21_input_sync_blk[3] | proc_21_output_sync_blk[3]);
    assign proc_21_data_FIFO_blk[4] = 1'b0;
    assign proc_21_data_PIPO_blk[4] = 1'b0;
    assign proc_21_start_FIFO_blk[4] = 1'b0;
    assign proc_21_TLF_FIFO_blk[4] = 1'b0;
    assign proc_21_input_sync_blk[4] = 1'b0;
    assign proc_21_output_sync_blk[4] = 1'b0 | (ap_done_reg_2 & write_back50_U0.ap_done & ~write_back51_U0.ap_done);
    assign proc_dep_vld_vec_21[4] = dl_detect_out ? proc_dep_vld_vec_21_reg[4] : (proc_21_data_FIFO_blk[4] | proc_21_data_PIPO_blk[4] | proc_21_start_FIFO_blk[4] | proc_21_TLF_FIFO_blk[4] | proc_21_input_sync_blk[4] | proc_21_output_sync_blk[4]);
    assign proc_21_data_FIFO_blk[5] = 1'b0;
    assign proc_21_data_PIPO_blk[5] = 1'b0;
    assign proc_21_start_FIFO_blk[5] = 1'b0;
    assign proc_21_TLF_FIFO_blk[5] = 1'b0;
    assign proc_21_input_sync_blk[5] = 1'b0;
    assign proc_21_output_sync_blk[5] = 1'b0 | (ap_done_reg_2 & write_back50_U0.ap_done & ~write_back52_U0.ap_done);
    assign proc_dep_vld_vec_21[5] = dl_detect_out ? proc_dep_vld_vec_21_reg[5] : (proc_21_data_FIFO_blk[5] | proc_21_data_PIPO_blk[5] | proc_21_start_FIFO_blk[5] | proc_21_TLF_FIFO_blk[5] | proc_21_input_sync_blk[5] | proc_21_output_sync_blk[5]);
    assign proc_21_data_FIFO_blk[6] = 1'b0;
    assign proc_21_data_PIPO_blk[6] = 1'b0;
    assign proc_21_start_FIFO_blk[6] = 1'b0;
    assign proc_21_TLF_FIFO_blk[6] = 1'b0;
    assign proc_21_input_sync_blk[6] = 1'b0;
    assign proc_21_output_sync_blk[6] = 1'b0 | (ap_done_reg_2 & write_back50_U0.ap_done & ~write_back53_U0.ap_done);
    assign proc_dep_vld_vec_21[6] = dl_detect_out ? proc_dep_vld_vec_21_reg[6] : (proc_21_data_FIFO_blk[6] | proc_21_data_PIPO_blk[6] | proc_21_start_FIFO_blk[6] | proc_21_TLF_FIFO_blk[6] | proc_21_input_sync_blk[6] | proc_21_output_sync_blk[6]);
    assign proc_21_data_FIFO_blk[7] = 1'b0;
    assign proc_21_data_PIPO_blk[7] = 1'b0;
    assign proc_21_start_FIFO_blk[7] = 1'b0;
    assign proc_21_TLF_FIFO_blk[7] = 1'b0;
    assign proc_21_input_sync_blk[7] = 1'b0;
    assign proc_21_output_sync_blk[7] = 1'b0 | (ap_done_reg_2 & write_back50_U0.ap_done & ~write_back54_U0.ap_done);
    assign proc_dep_vld_vec_21[7] = dl_detect_out ? proc_dep_vld_vec_21_reg[7] : (proc_21_data_FIFO_blk[7] | proc_21_data_PIPO_blk[7] | proc_21_start_FIFO_blk[7] | proc_21_TLF_FIFO_blk[7] | proc_21_input_sync_blk[7] | proc_21_output_sync_blk[7]);
    assign proc_21_data_FIFO_blk[8] = 1'b0;
    assign proc_21_data_PIPO_blk[8] = 1'b0;
    assign proc_21_start_FIFO_blk[8] = 1'b0;
    assign proc_21_TLF_FIFO_blk[8] = 1'b0;
    assign proc_21_input_sync_blk[8] = 1'b0;
    assign proc_21_output_sync_blk[8] = 1'b0 | (ap_done_reg_2 & write_back50_U0.ap_done & ~write_back55_U0.ap_done);
    assign proc_dep_vld_vec_21[8] = dl_detect_out ? proc_dep_vld_vec_21_reg[8] : (proc_21_data_FIFO_blk[8] | proc_21_data_PIPO_blk[8] | proc_21_start_FIFO_blk[8] | proc_21_TLF_FIFO_blk[8] | proc_21_input_sync_blk[8] | proc_21_output_sync_blk[8]);
    assign proc_21_data_FIFO_blk[9] = 1'b0;
    assign proc_21_data_PIPO_blk[9] = 1'b0;
    assign proc_21_start_FIFO_blk[9] = 1'b0;
    assign proc_21_TLF_FIFO_blk[9] = 1'b0;
    assign proc_21_input_sync_blk[9] = 1'b0;
    assign proc_21_output_sync_blk[9] = 1'b0 | (ap_done_reg_2 & write_back50_U0.ap_done & ~write_back56_U0.ap_done);
    assign proc_dep_vld_vec_21[9] = dl_detect_out ? proc_dep_vld_vec_21_reg[9] : (proc_21_data_FIFO_blk[9] | proc_21_data_PIPO_blk[9] | proc_21_start_FIFO_blk[9] | proc_21_TLF_FIFO_blk[9] | proc_21_input_sync_blk[9] | proc_21_output_sync_blk[9]);
    assign proc_21_data_FIFO_blk[10] = 1'b0;
    assign proc_21_data_PIPO_blk[10] = 1'b0;
    assign proc_21_start_FIFO_blk[10] = 1'b0;
    assign proc_21_TLF_FIFO_blk[10] = 1'b0;
    assign proc_21_input_sync_blk[10] = 1'b0;
    assign proc_21_output_sync_blk[10] = 1'b0 | (ap_done_reg_2 & write_back50_U0.ap_done & ~write_back57_U0.ap_done);
    assign proc_dep_vld_vec_21[10] = dl_detect_out ? proc_dep_vld_vec_21_reg[10] : (proc_21_data_FIFO_blk[10] | proc_21_data_PIPO_blk[10] | proc_21_start_FIFO_blk[10] | proc_21_TLF_FIFO_blk[10] | proc_21_input_sync_blk[10] | proc_21_output_sync_blk[10]);
    assign proc_21_data_FIFO_blk[11] = 1'b0;
    assign proc_21_data_PIPO_blk[11] = 1'b0;
    assign proc_21_start_FIFO_blk[11] = 1'b0;
    assign proc_21_TLF_FIFO_blk[11] = 1'b0;
    assign proc_21_input_sync_blk[11] = 1'b0;
    assign proc_21_output_sync_blk[11] = 1'b0 | (ap_done_reg_2 & write_back50_U0.ap_done & ~write_back58_U0.ap_done);
    assign proc_dep_vld_vec_21[11] = dl_detect_out ? proc_dep_vld_vec_21_reg[11] : (proc_21_data_FIFO_blk[11] | proc_21_data_PIPO_blk[11] | proc_21_start_FIFO_blk[11] | proc_21_TLF_FIFO_blk[11] | proc_21_input_sync_blk[11] | proc_21_output_sync_blk[11]);
    assign proc_21_data_FIFO_blk[12] = 1'b0;
    assign proc_21_data_PIPO_blk[12] = 1'b0;
    assign proc_21_start_FIFO_blk[12] = 1'b0;
    assign proc_21_TLF_FIFO_blk[12] = 1'b0;
    assign proc_21_input_sync_blk[12] = 1'b0;
    assign proc_21_output_sync_blk[12] = 1'b0 | (ap_done_reg_2 & write_back50_U0.ap_done & ~write_back59_U0.ap_done);
    assign proc_dep_vld_vec_21[12] = dl_detect_out ? proc_dep_vld_vec_21_reg[12] : (proc_21_data_FIFO_blk[12] | proc_21_data_PIPO_blk[12] | proc_21_start_FIFO_blk[12] | proc_21_TLF_FIFO_blk[12] | proc_21_input_sync_blk[12] | proc_21_output_sync_blk[12]);
    assign proc_21_data_FIFO_blk[13] = 1'b0;
    assign proc_21_data_PIPO_blk[13] = 1'b0;
    assign proc_21_start_FIFO_blk[13] = 1'b0;
    assign proc_21_TLF_FIFO_blk[13] = 1'b0;
    assign proc_21_input_sync_blk[13] = 1'b0;
    assign proc_21_output_sync_blk[13] = 1'b0 | (ap_done_reg_2 & write_back50_U0.ap_done & ~write_back60_U0.ap_done);
    assign proc_dep_vld_vec_21[13] = dl_detect_out ? proc_dep_vld_vec_21_reg[13] : (proc_21_data_FIFO_blk[13] | proc_21_data_PIPO_blk[13] | proc_21_start_FIFO_blk[13] | proc_21_TLF_FIFO_blk[13] | proc_21_input_sync_blk[13] | proc_21_output_sync_blk[13]);
    assign proc_21_data_FIFO_blk[14] = 1'b0;
    assign proc_21_data_PIPO_blk[14] = 1'b0;
    assign proc_21_start_FIFO_blk[14] = 1'b0;
    assign proc_21_TLF_FIFO_blk[14] = 1'b0;
    assign proc_21_input_sync_blk[14] = 1'b0;
    assign proc_21_output_sync_blk[14] = 1'b0 | (ap_done_reg_2 & write_back50_U0.ap_done & ~write_back61_U0.ap_done);
    assign proc_dep_vld_vec_21[14] = dl_detect_out ? proc_dep_vld_vec_21_reg[14] : (proc_21_data_FIFO_blk[14] | proc_21_data_PIPO_blk[14] | proc_21_start_FIFO_blk[14] | proc_21_TLF_FIFO_blk[14] | proc_21_input_sync_blk[14] | proc_21_output_sync_blk[14]);
    assign proc_21_data_FIFO_blk[15] = 1'b0;
    assign proc_21_data_PIPO_blk[15] = 1'b0;
    assign proc_21_start_FIFO_blk[15] = 1'b0;
    assign proc_21_TLF_FIFO_blk[15] = 1'b0;
    assign proc_21_input_sync_blk[15] = 1'b0;
    assign proc_21_output_sync_blk[15] = 1'b0 | (ap_done_reg_2 & write_back50_U0.ap_done & ~write_back62_U0.ap_done);
    assign proc_dep_vld_vec_21[15] = dl_detect_out ? proc_dep_vld_vec_21_reg[15] : (proc_21_data_FIFO_blk[15] | proc_21_data_PIPO_blk[15] | proc_21_start_FIFO_blk[15] | proc_21_TLF_FIFO_blk[15] | proc_21_input_sync_blk[15] | proc_21_output_sync_blk[15]);
    assign proc_21_data_FIFO_blk[16] = 1'b0;
    assign proc_21_data_PIPO_blk[16] = 1'b0;
    assign proc_21_start_FIFO_blk[16] = 1'b0;
    assign proc_21_TLF_FIFO_blk[16] = 1'b0;
    assign proc_21_input_sync_blk[16] = 1'b0;
    assign proc_21_output_sync_blk[16] = 1'b0 | (ap_done_reg_2 & write_back50_U0.ap_done & ~write_back63_U0.ap_done);
    assign proc_dep_vld_vec_21[16] = dl_detect_out ? proc_dep_vld_vec_21_reg[16] : (proc_21_data_FIFO_blk[16] | proc_21_data_PIPO_blk[16] | proc_21_start_FIFO_blk[16] | proc_21_TLF_FIFO_blk[16] | proc_21_input_sync_blk[16] | proc_21_output_sync_blk[16]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_21_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_21_reg <= proc_dep_vld_vec_21;
        end
    end
    assign in_chan_dep_vld_vec_21[0] = dep_chan_vld_0_21;
    assign in_chan_dep_data_vec_21[34 : 0] = dep_chan_data_0_21;
    assign token_in_vec_21[0] = token_0_21;
    assign in_chan_dep_vld_vec_21[1] = dep_chan_vld_5_21;
    assign in_chan_dep_data_vec_21[69 : 35] = dep_chan_data_5_21;
    assign token_in_vec_21[1] = token_5_21;
    assign in_chan_dep_vld_vec_21[2] = dep_chan_vld_19_21;
    assign in_chan_dep_data_vec_21[104 : 70] = dep_chan_data_19_21;
    assign token_in_vec_21[2] = token_19_21;
    assign in_chan_dep_vld_vec_21[3] = dep_chan_vld_20_21;
    assign in_chan_dep_data_vec_21[139 : 105] = dep_chan_data_20_21;
    assign token_in_vec_21[3] = token_20_21;
    assign in_chan_dep_vld_vec_21[4] = dep_chan_vld_22_21;
    assign in_chan_dep_data_vec_21[174 : 140] = dep_chan_data_22_21;
    assign token_in_vec_21[4] = token_22_21;
    assign in_chan_dep_vld_vec_21[5] = dep_chan_vld_23_21;
    assign in_chan_dep_data_vec_21[209 : 175] = dep_chan_data_23_21;
    assign token_in_vec_21[5] = token_23_21;
    assign in_chan_dep_vld_vec_21[6] = dep_chan_vld_24_21;
    assign in_chan_dep_data_vec_21[244 : 210] = dep_chan_data_24_21;
    assign token_in_vec_21[6] = token_24_21;
    assign in_chan_dep_vld_vec_21[7] = dep_chan_vld_25_21;
    assign in_chan_dep_data_vec_21[279 : 245] = dep_chan_data_25_21;
    assign token_in_vec_21[7] = token_25_21;
    assign in_chan_dep_vld_vec_21[8] = dep_chan_vld_26_21;
    assign in_chan_dep_data_vec_21[314 : 280] = dep_chan_data_26_21;
    assign token_in_vec_21[8] = token_26_21;
    assign in_chan_dep_vld_vec_21[9] = dep_chan_vld_27_21;
    assign in_chan_dep_data_vec_21[349 : 315] = dep_chan_data_27_21;
    assign token_in_vec_21[9] = token_27_21;
    assign in_chan_dep_vld_vec_21[10] = dep_chan_vld_28_21;
    assign in_chan_dep_data_vec_21[384 : 350] = dep_chan_data_28_21;
    assign token_in_vec_21[10] = token_28_21;
    assign in_chan_dep_vld_vec_21[11] = dep_chan_vld_29_21;
    assign in_chan_dep_data_vec_21[419 : 385] = dep_chan_data_29_21;
    assign token_in_vec_21[11] = token_29_21;
    assign in_chan_dep_vld_vec_21[12] = dep_chan_vld_30_21;
    assign in_chan_dep_data_vec_21[454 : 420] = dep_chan_data_30_21;
    assign token_in_vec_21[12] = token_30_21;
    assign in_chan_dep_vld_vec_21[13] = dep_chan_vld_31_21;
    assign in_chan_dep_data_vec_21[489 : 455] = dep_chan_data_31_21;
    assign token_in_vec_21[13] = token_31_21;
    assign in_chan_dep_vld_vec_21[14] = dep_chan_vld_32_21;
    assign in_chan_dep_data_vec_21[524 : 490] = dep_chan_data_32_21;
    assign token_in_vec_21[14] = token_32_21;
    assign in_chan_dep_vld_vec_21[15] = dep_chan_vld_33_21;
    assign in_chan_dep_data_vec_21[559 : 525] = dep_chan_data_33_21;
    assign token_in_vec_21[15] = token_33_21;
    assign in_chan_dep_vld_vec_21[16] = dep_chan_vld_34_21;
    assign in_chan_dep_data_vec_21[594 : 560] = dep_chan_data_34_21;
    assign token_in_vec_21[16] = token_34_21;
    assign dep_chan_vld_21_0 = out_chan_dep_vld_vec_21[0];
    assign dep_chan_data_21_0 = out_chan_dep_data_21;
    assign token_21_0 = token_out_vec_21[0];
    assign dep_chan_vld_21_5 = out_chan_dep_vld_vec_21[1];
    assign dep_chan_data_21_5 = out_chan_dep_data_21;
    assign token_21_5 = token_out_vec_21[1];
    assign dep_chan_vld_21_19 = out_chan_dep_vld_vec_21[2];
    assign dep_chan_data_21_19 = out_chan_dep_data_21;
    assign token_21_19 = token_out_vec_21[2];
    assign dep_chan_vld_21_20 = out_chan_dep_vld_vec_21[3];
    assign dep_chan_data_21_20 = out_chan_dep_data_21;
    assign token_21_20 = token_out_vec_21[3];
    assign dep_chan_vld_21_22 = out_chan_dep_vld_vec_21[4];
    assign dep_chan_data_21_22 = out_chan_dep_data_21;
    assign token_21_22 = token_out_vec_21[4];
    assign dep_chan_vld_21_23 = out_chan_dep_vld_vec_21[5];
    assign dep_chan_data_21_23 = out_chan_dep_data_21;
    assign token_21_23 = token_out_vec_21[5];
    assign dep_chan_vld_21_24 = out_chan_dep_vld_vec_21[6];
    assign dep_chan_data_21_24 = out_chan_dep_data_21;
    assign token_21_24 = token_out_vec_21[6];
    assign dep_chan_vld_21_25 = out_chan_dep_vld_vec_21[7];
    assign dep_chan_data_21_25 = out_chan_dep_data_21;
    assign token_21_25 = token_out_vec_21[7];
    assign dep_chan_vld_21_26 = out_chan_dep_vld_vec_21[8];
    assign dep_chan_data_21_26 = out_chan_dep_data_21;
    assign token_21_26 = token_out_vec_21[8];
    assign dep_chan_vld_21_27 = out_chan_dep_vld_vec_21[9];
    assign dep_chan_data_21_27 = out_chan_dep_data_21;
    assign token_21_27 = token_out_vec_21[9];
    assign dep_chan_vld_21_28 = out_chan_dep_vld_vec_21[10];
    assign dep_chan_data_21_28 = out_chan_dep_data_21;
    assign token_21_28 = token_out_vec_21[10];
    assign dep_chan_vld_21_29 = out_chan_dep_vld_vec_21[11];
    assign dep_chan_data_21_29 = out_chan_dep_data_21;
    assign token_21_29 = token_out_vec_21[11];
    assign dep_chan_vld_21_30 = out_chan_dep_vld_vec_21[12];
    assign dep_chan_data_21_30 = out_chan_dep_data_21;
    assign token_21_30 = token_out_vec_21[12];
    assign dep_chan_vld_21_31 = out_chan_dep_vld_vec_21[13];
    assign dep_chan_data_21_31 = out_chan_dep_data_21;
    assign token_21_31 = token_out_vec_21[13];
    assign dep_chan_vld_21_32 = out_chan_dep_vld_vec_21[14];
    assign dep_chan_data_21_32 = out_chan_dep_data_21;
    assign token_21_32 = token_out_vec_21[14];
    assign dep_chan_vld_21_33 = out_chan_dep_vld_vec_21[15];
    assign dep_chan_data_21_33 = out_chan_dep_data_21;
    assign token_21_33 = token_out_vec_21[15];
    assign dep_chan_vld_21_34 = out_chan_dep_vld_vec_21[16];
    assign dep_chan_data_21_34 = out_chan_dep_data_21;
    assign token_21_34 = token_out_vec_21[16];

    // Process: write_back51_U0
    kernel_pr_hls_deadlock_detect_unit #(35, 22, 17, 17) kernel_pr_hls_deadlock_detect_unit_22 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_22),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_22),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_22),
        .token_in_vec(token_in_vec_22),
        .dl_detect_in(dl_detect_out),
        .origin(origin[22]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_22),
        .out_chan_dep_data(out_chan_dep_data_22),
        .token_out_vec(token_out_vec_22),
        .dl_detect_out(dl_in_vec[22]));

    assign proc_22_data_FIFO_blk[0] = 1'b0 | (~write_back51_U0.H_blk_n) | (~write_back51_U0.hyperedge_size_blk_n);
    assign proc_22_data_PIPO_blk[0] = 1'b0;
    assign proc_22_start_FIFO_blk[0] = 1'b0 | (~start_for_write_back51_U0_U.if_empty_n & write_back51_U0.ap_idle & ~start_for_write_back51_U0_U.if_write);
    assign proc_22_TLF_FIFO_blk[0] = 1'b0;
    assign proc_22_input_sync_blk[0] = 1'b0;
    assign proc_22_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_22[0] = dl_detect_out ? proc_dep_vld_vec_22_reg[0] : (proc_22_data_FIFO_blk[0] | proc_22_data_PIPO_blk[0] | proc_22_start_FIFO_blk[0] | proc_22_TLF_FIFO_blk[0] | proc_22_input_sync_blk[0] | proc_22_output_sync_blk[0]);
    assign proc_22_data_FIFO_blk[1] = 1'b0 | (~write_back51_U0.value_stream_V_V3_blk_n);
    assign proc_22_data_PIPO_blk[1] = 1'b0;
    assign proc_22_start_FIFO_blk[1] = 1'b0;
    assign proc_22_TLF_FIFO_blk[1] = 1'b0;
    assign proc_22_input_sync_blk[1] = 1'b0;
    assign proc_22_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_22[1] = dl_detect_out ? proc_dep_vld_vec_22_reg[1] : (proc_22_data_FIFO_blk[1] | proc_22_data_PIPO_blk[1] | proc_22_start_FIFO_blk[1] | proc_22_TLF_FIFO_blk[1] | proc_22_input_sync_blk[1] | proc_22_output_sync_blk[1]);
    assign proc_22_data_FIFO_blk[2] = 1'b0;
    assign proc_22_data_PIPO_blk[2] = 1'b0;
    assign proc_22_start_FIFO_blk[2] = 1'b0;
    assign proc_22_TLF_FIFO_blk[2] = 1'b0;
    assign proc_22_input_sync_blk[2] = 1'b0;
    assign proc_22_output_sync_blk[2] = 1'b0 | (ap_done_reg_3 & write_back51_U0.ap_done & ~write_back48_U0.ap_done);
    assign proc_dep_vld_vec_22[2] = dl_detect_out ? proc_dep_vld_vec_22_reg[2] : (proc_22_data_FIFO_blk[2] | proc_22_data_PIPO_blk[2] | proc_22_start_FIFO_blk[2] | proc_22_TLF_FIFO_blk[2] | proc_22_input_sync_blk[2] | proc_22_output_sync_blk[2]);
    assign proc_22_data_FIFO_blk[3] = 1'b0;
    assign proc_22_data_PIPO_blk[3] = 1'b0;
    assign proc_22_start_FIFO_blk[3] = 1'b0;
    assign proc_22_TLF_FIFO_blk[3] = 1'b0;
    assign proc_22_input_sync_blk[3] = 1'b0;
    assign proc_22_output_sync_blk[3] = 1'b0 | (ap_done_reg_3 & write_back51_U0.ap_done & ~write_back49_U0.ap_done);
    assign proc_dep_vld_vec_22[3] = dl_detect_out ? proc_dep_vld_vec_22_reg[3] : (proc_22_data_FIFO_blk[3] | proc_22_data_PIPO_blk[3] | proc_22_start_FIFO_blk[3] | proc_22_TLF_FIFO_blk[3] | proc_22_input_sync_blk[3] | proc_22_output_sync_blk[3]);
    assign proc_22_data_FIFO_blk[4] = 1'b0;
    assign proc_22_data_PIPO_blk[4] = 1'b0;
    assign proc_22_start_FIFO_blk[4] = 1'b0;
    assign proc_22_TLF_FIFO_blk[4] = 1'b0;
    assign proc_22_input_sync_blk[4] = 1'b0;
    assign proc_22_output_sync_blk[4] = 1'b0 | (ap_done_reg_3 & write_back51_U0.ap_done & ~write_back50_U0.ap_done);
    assign proc_dep_vld_vec_22[4] = dl_detect_out ? proc_dep_vld_vec_22_reg[4] : (proc_22_data_FIFO_blk[4] | proc_22_data_PIPO_blk[4] | proc_22_start_FIFO_blk[4] | proc_22_TLF_FIFO_blk[4] | proc_22_input_sync_blk[4] | proc_22_output_sync_blk[4]);
    assign proc_22_data_FIFO_blk[5] = 1'b0;
    assign proc_22_data_PIPO_blk[5] = 1'b0;
    assign proc_22_start_FIFO_blk[5] = 1'b0;
    assign proc_22_TLF_FIFO_blk[5] = 1'b0;
    assign proc_22_input_sync_blk[5] = 1'b0;
    assign proc_22_output_sync_blk[5] = 1'b0 | (ap_done_reg_3 & write_back51_U0.ap_done & ~write_back52_U0.ap_done);
    assign proc_dep_vld_vec_22[5] = dl_detect_out ? proc_dep_vld_vec_22_reg[5] : (proc_22_data_FIFO_blk[5] | proc_22_data_PIPO_blk[5] | proc_22_start_FIFO_blk[5] | proc_22_TLF_FIFO_blk[5] | proc_22_input_sync_blk[5] | proc_22_output_sync_blk[5]);
    assign proc_22_data_FIFO_blk[6] = 1'b0;
    assign proc_22_data_PIPO_blk[6] = 1'b0;
    assign proc_22_start_FIFO_blk[6] = 1'b0;
    assign proc_22_TLF_FIFO_blk[6] = 1'b0;
    assign proc_22_input_sync_blk[6] = 1'b0;
    assign proc_22_output_sync_blk[6] = 1'b0 | (ap_done_reg_3 & write_back51_U0.ap_done & ~write_back53_U0.ap_done);
    assign proc_dep_vld_vec_22[6] = dl_detect_out ? proc_dep_vld_vec_22_reg[6] : (proc_22_data_FIFO_blk[6] | proc_22_data_PIPO_blk[6] | proc_22_start_FIFO_blk[6] | proc_22_TLF_FIFO_blk[6] | proc_22_input_sync_blk[6] | proc_22_output_sync_blk[6]);
    assign proc_22_data_FIFO_blk[7] = 1'b0;
    assign proc_22_data_PIPO_blk[7] = 1'b0;
    assign proc_22_start_FIFO_blk[7] = 1'b0;
    assign proc_22_TLF_FIFO_blk[7] = 1'b0;
    assign proc_22_input_sync_blk[7] = 1'b0;
    assign proc_22_output_sync_blk[7] = 1'b0 | (ap_done_reg_3 & write_back51_U0.ap_done & ~write_back54_U0.ap_done);
    assign proc_dep_vld_vec_22[7] = dl_detect_out ? proc_dep_vld_vec_22_reg[7] : (proc_22_data_FIFO_blk[7] | proc_22_data_PIPO_blk[7] | proc_22_start_FIFO_blk[7] | proc_22_TLF_FIFO_blk[7] | proc_22_input_sync_blk[7] | proc_22_output_sync_blk[7]);
    assign proc_22_data_FIFO_blk[8] = 1'b0;
    assign proc_22_data_PIPO_blk[8] = 1'b0;
    assign proc_22_start_FIFO_blk[8] = 1'b0;
    assign proc_22_TLF_FIFO_blk[8] = 1'b0;
    assign proc_22_input_sync_blk[8] = 1'b0;
    assign proc_22_output_sync_blk[8] = 1'b0 | (ap_done_reg_3 & write_back51_U0.ap_done & ~write_back55_U0.ap_done);
    assign proc_dep_vld_vec_22[8] = dl_detect_out ? proc_dep_vld_vec_22_reg[8] : (proc_22_data_FIFO_blk[8] | proc_22_data_PIPO_blk[8] | proc_22_start_FIFO_blk[8] | proc_22_TLF_FIFO_blk[8] | proc_22_input_sync_blk[8] | proc_22_output_sync_blk[8]);
    assign proc_22_data_FIFO_blk[9] = 1'b0;
    assign proc_22_data_PIPO_blk[9] = 1'b0;
    assign proc_22_start_FIFO_blk[9] = 1'b0;
    assign proc_22_TLF_FIFO_blk[9] = 1'b0;
    assign proc_22_input_sync_blk[9] = 1'b0;
    assign proc_22_output_sync_blk[9] = 1'b0 | (ap_done_reg_3 & write_back51_U0.ap_done & ~write_back56_U0.ap_done);
    assign proc_dep_vld_vec_22[9] = dl_detect_out ? proc_dep_vld_vec_22_reg[9] : (proc_22_data_FIFO_blk[9] | proc_22_data_PIPO_blk[9] | proc_22_start_FIFO_blk[9] | proc_22_TLF_FIFO_blk[9] | proc_22_input_sync_blk[9] | proc_22_output_sync_blk[9]);
    assign proc_22_data_FIFO_blk[10] = 1'b0;
    assign proc_22_data_PIPO_blk[10] = 1'b0;
    assign proc_22_start_FIFO_blk[10] = 1'b0;
    assign proc_22_TLF_FIFO_blk[10] = 1'b0;
    assign proc_22_input_sync_blk[10] = 1'b0;
    assign proc_22_output_sync_blk[10] = 1'b0 | (ap_done_reg_3 & write_back51_U0.ap_done & ~write_back57_U0.ap_done);
    assign proc_dep_vld_vec_22[10] = dl_detect_out ? proc_dep_vld_vec_22_reg[10] : (proc_22_data_FIFO_blk[10] | proc_22_data_PIPO_blk[10] | proc_22_start_FIFO_blk[10] | proc_22_TLF_FIFO_blk[10] | proc_22_input_sync_blk[10] | proc_22_output_sync_blk[10]);
    assign proc_22_data_FIFO_blk[11] = 1'b0;
    assign proc_22_data_PIPO_blk[11] = 1'b0;
    assign proc_22_start_FIFO_blk[11] = 1'b0;
    assign proc_22_TLF_FIFO_blk[11] = 1'b0;
    assign proc_22_input_sync_blk[11] = 1'b0;
    assign proc_22_output_sync_blk[11] = 1'b0 | (ap_done_reg_3 & write_back51_U0.ap_done & ~write_back58_U0.ap_done);
    assign proc_dep_vld_vec_22[11] = dl_detect_out ? proc_dep_vld_vec_22_reg[11] : (proc_22_data_FIFO_blk[11] | proc_22_data_PIPO_blk[11] | proc_22_start_FIFO_blk[11] | proc_22_TLF_FIFO_blk[11] | proc_22_input_sync_blk[11] | proc_22_output_sync_blk[11]);
    assign proc_22_data_FIFO_blk[12] = 1'b0;
    assign proc_22_data_PIPO_blk[12] = 1'b0;
    assign proc_22_start_FIFO_blk[12] = 1'b0;
    assign proc_22_TLF_FIFO_blk[12] = 1'b0;
    assign proc_22_input_sync_blk[12] = 1'b0;
    assign proc_22_output_sync_blk[12] = 1'b0 | (ap_done_reg_3 & write_back51_U0.ap_done & ~write_back59_U0.ap_done);
    assign proc_dep_vld_vec_22[12] = dl_detect_out ? proc_dep_vld_vec_22_reg[12] : (proc_22_data_FIFO_blk[12] | proc_22_data_PIPO_blk[12] | proc_22_start_FIFO_blk[12] | proc_22_TLF_FIFO_blk[12] | proc_22_input_sync_blk[12] | proc_22_output_sync_blk[12]);
    assign proc_22_data_FIFO_blk[13] = 1'b0;
    assign proc_22_data_PIPO_blk[13] = 1'b0;
    assign proc_22_start_FIFO_blk[13] = 1'b0;
    assign proc_22_TLF_FIFO_blk[13] = 1'b0;
    assign proc_22_input_sync_blk[13] = 1'b0;
    assign proc_22_output_sync_blk[13] = 1'b0 | (ap_done_reg_3 & write_back51_U0.ap_done & ~write_back60_U0.ap_done);
    assign proc_dep_vld_vec_22[13] = dl_detect_out ? proc_dep_vld_vec_22_reg[13] : (proc_22_data_FIFO_blk[13] | proc_22_data_PIPO_blk[13] | proc_22_start_FIFO_blk[13] | proc_22_TLF_FIFO_blk[13] | proc_22_input_sync_blk[13] | proc_22_output_sync_blk[13]);
    assign proc_22_data_FIFO_blk[14] = 1'b0;
    assign proc_22_data_PIPO_blk[14] = 1'b0;
    assign proc_22_start_FIFO_blk[14] = 1'b0;
    assign proc_22_TLF_FIFO_blk[14] = 1'b0;
    assign proc_22_input_sync_blk[14] = 1'b0;
    assign proc_22_output_sync_blk[14] = 1'b0 | (ap_done_reg_3 & write_back51_U0.ap_done & ~write_back61_U0.ap_done);
    assign proc_dep_vld_vec_22[14] = dl_detect_out ? proc_dep_vld_vec_22_reg[14] : (proc_22_data_FIFO_blk[14] | proc_22_data_PIPO_blk[14] | proc_22_start_FIFO_blk[14] | proc_22_TLF_FIFO_blk[14] | proc_22_input_sync_blk[14] | proc_22_output_sync_blk[14]);
    assign proc_22_data_FIFO_blk[15] = 1'b0;
    assign proc_22_data_PIPO_blk[15] = 1'b0;
    assign proc_22_start_FIFO_blk[15] = 1'b0;
    assign proc_22_TLF_FIFO_blk[15] = 1'b0;
    assign proc_22_input_sync_blk[15] = 1'b0;
    assign proc_22_output_sync_blk[15] = 1'b0 | (ap_done_reg_3 & write_back51_U0.ap_done & ~write_back62_U0.ap_done);
    assign proc_dep_vld_vec_22[15] = dl_detect_out ? proc_dep_vld_vec_22_reg[15] : (proc_22_data_FIFO_blk[15] | proc_22_data_PIPO_blk[15] | proc_22_start_FIFO_blk[15] | proc_22_TLF_FIFO_blk[15] | proc_22_input_sync_blk[15] | proc_22_output_sync_blk[15]);
    assign proc_22_data_FIFO_blk[16] = 1'b0;
    assign proc_22_data_PIPO_blk[16] = 1'b0;
    assign proc_22_start_FIFO_blk[16] = 1'b0;
    assign proc_22_TLF_FIFO_blk[16] = 1'b0;
    assign proc_22_input_sync_blk[16] = 1'b0;
    assign proc_22_output_sync_blk[16] = 1'b0 | (ap_done_reg_3 & write_back51_U0.ap_done & ~write_back63_U0.ap_done);
    assign proc_dep_vld_vec_22[16] = dl_detect_out ? proc_dep_vld_vec_22_reg[16] : (proc_22_data_FIFO_blk[16] | proc_22_data_PIPO_blk[16] | proc_22_start_FIFO_blk[16] | proc_22_TLF_FIFO_blk[16] | proc_22_input_sync_blk[16] | proc_22_output_sync_blk[16]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_22_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_22_reg <= proc_dep_vld_vec_22;
        end
    end
    assign in_chan_dep_vld_vec_22[0] = dep_chan_vld_0_22;
    assign in_chan_dep_data_vec_22[34 : 0] = dep_chan_data_0_22;
    assign token_in_vec_22[0] = token_0_22;
    assign in_chan_dep_vld_vec_22[1] = dep_chan_vld_6_22;
    assign in_chan_dep_data_vec_22[69 : 35] = dep_chan_data_6_22;
    assign token_in_vec_22[1] = token_6_22;
    assign in_chan_dep_vld_vec_22[2] = dep_chan_vld_19_22;
    assign in_chan_dep_data_vec_22[104 : 70] = dep_chan_data_19_22;
    assign token_in_vec_22[2] = token_19_22;
    assign in_chan_dep_vld_vec_22[3] = dep_chan_vld_20_22;
    assign in_chan_dep_data_vec_22[139 : 105] = dep_chan_data_20_22;
    assign token_in_vec_22[3] = token_20_22;
    assign in_chan_dep_vld_vec_22[4] = dep_chan_vld_21_22;
    assign in_chan_dep_data_vec_22[174 : 140] = dep_chan_data_21_22;
    assign token_in_vec_22[4] = token_21_22;
    assign in_chan_dep_vld_vec_22[5] = dep_chan_vld_23_22;
    assign in_chan_dep_data_vec_22[209 : 175] = dep_chan_data_23_22;
    assign token_in_vec_22[5] = token_23_22;
    assign in_chan_dep_vld_vec_22[6] = dep_chan_vld_24_22;
    assign in_chan_dep_data_vec_22[244 : 210] = dep_chan_data_24_22;
    assign token_in_vec_22[6] = token_24_22;
    assign in_chan_dep_vld_vec_22[7] = dep_chan_vld_25_22;
    assign in_chan_dep_data_vec_22[279 : 245] = dep_chan_data_25_22;
    assign token_in_vec_22[7] = token_25_22;
    assign in_chan_dep_vld_vec_22[8] = dep_chan_vld_26_22;
    assign in_chan_dep_data_vec_22[314 : 280] = dep_chan_data_26_22;
    assign token_in_vec_22[8] = token_26_22;
    assign in_chan_dep_vld_vec_22[9] = dep_chan_vld_27_22;
    assign in_chan_dep_data_vec_22[349 : 315] = dep_chan_data_27_22;
    assign token_in_vec_22[9] = token_27_22;
    assign in_chan_dep_vld_vec_22[10] = dep_chan_vld_28_22;
    assign in_chan_dep_data_vec_22[384 : 350] = dep_chan_data_28_22;
    assign token_in_vec_22[10] = token_28_22;
    assign in_chan_dep_vld_vec_22[11] = dep_chan_vld_29_22;
    assign in_chan_dep_data_vec_22[419 : 385] = dep_chan_data_29_22;
    assign token_in_vec_22[11] = token_29_22;
    assign in_chan_dep_vld_vec_22[12] = dep_chan_vld_30_22;
    assign in_chan_dep_data_vec_22[454 : 420] = dep_chan_data_30_22;
    assign token_in_vec_22[12] = token_30_22;
    assign in_chan_dep_vld_vec_22[13] = dep_chan_vld_31_22;
    assign in_chan_dep_data_vec_22[489 : 455] = dep_chan_data_31_22;
    assign token_in_vec_22[13] = token_31_22;
    assign in_chan_dep_vld_vec_22[14] = dep_chan_vld_32_22;
    assign in_chan_dep_data_vec_22[524 : 490] = dep_chan_data_32_22;
    assign token_in_vec_22[14] = token_32_22;
    assign in_chan_dep_vld_vec_22[15] = dep_chan_vld_33_22;
    assign in_chan_dep_data_vec_22[559 : 525] = dep_chan_data_33_22;
    assign token_in_vec_22[15] = token_33_22;
    assign in_chan_dep_vld_vec_22[16] = dep_chan_vld_34_22;
    assign in_chan_dep_data_vec_22[594 : 560] = dep_chan_data_34_22;
    assign token_in_vec_22[16] = token_34_22;
    assign dep_chan_vld_22_0 = out_chan_dep_vld_vec_22[0];
    assign dep_chan_data_22_0 = out_chan_dep_data_22;
    assign token_22_0 = token_out_vec_22[0];
    assign dep_chan_vld_22_6 = out_chan_dep_vld_vec_22[1];
    assign dep_chan_data_22_6 = out_chan_dep_data_22;
    assign token_22_6 = token_out_vec_22[1];
    assign dep_chan_vld_22_19 = out_chan_dep_vld_vec_22[2];
    assign dep_chan_data_22_19 = out_chan_dep_data_22;
    assign token_22_19 = token_out_vec_22[2];
    assign dep_chan_vld_22_20 = out_chan_dep_vld_vec_22[3];
    assign dep_chan_data_22_20 = out_chan_dep_data_22;
    assign token_22_20 = token_out_vec_22[3];
    assign dep_chan_vld_22_21 = out_chan_dep_vld_vec_22[4];
    assign dep_chan_data_22_21 = out_chan_dep_data_22;
    assign token_22_21 = token_out_vec_22[4];
    assign dep_chan_vld_22_23 = out_chan_dep_vld_vec_22[5];
    assign dep_chan_data_22_23 = out_chan_dep_data_22;
    assign token_22_23 = token_out_vec_22[5];
    assign dep_chan_vld_22_24 = out_chan_dep_vld_vec_22[6];
    assign dep_chan_data_22_24 = out_chan_dep_data_22;
    assign token_22_24 = token_out_vec_22[6];
    assign dep_chan_vld_22_25 = out_chan_dep_vld_vec_22[7];
    assign dep_chan_data_22_25 = out_chan_dep_data_22;
    assign token_22_25 = token_out_vec_22[7];
    assign dep_chan_vld_22_26 = out_chan_dep_vld_vec_22[8];
    assign dep_chan_data_22_26 = out_chan_dep_data_22;
    assign token_22_26 = token_out_vec_22[8];
    assign dep_chan_vld_22_27 = out_chan_dep_vld_vec_22[9];
    assign dep_chan_data_22_27 = out_chan_dep_data_22;
    assign token_22_27 = token_out_vec_22[9];
    assign dep_chan_vld_22_28 = out_chan_dep_vld_vec_22[10];
    assign dep_chan_data_22_28 = out_chan_dep_data_22;
    assign token_22_28 = token_out_vec_22[10];
    assign dep_chan_vld_22_29 = out_chan_dep_vld_vec_22[11];
    assign dep_chan_data_22_29 = out_chan_dep_data_22;
    assign token_22_29 = token_out_vec_22[11];
    assign dep_chan_vld_22_30 = out_chan_dep_vld_vec_22[12];
    assign dep_chan_data_22_30 = out_chan_dep_data_22;
    assign token_22_30 = token_out_vec_22[12];
    assign dep_chan_vld_22_31 = out_chan_dep_vld_vec_22[13];
    assign dep_chan_data_22_31 = out_chan_dep_data_22;
    assign token_22_31 = token_out_vec_22[13];
    assign dep_chan_vld_22_32 = out_chan_dep_vld_vec_22[14];
    assign dep_chan_data_22_32 = out_chan_dep_data_22;
    assign token_22_32 = token_out_vec_22[14];
    assign dep_chan_vld_22_33 = out_chan_dep_vld_vec_22[15];
    assign dep_chan_data_22_33 = out_chan_dep_data_22;
    assign token_22_33 = token_out_vec_22[15];
    assign dep_chan_vld_22_34 = out_chan_dep_vld_vec_22[16];
    assign dep_chan_data_22_34 = out_chan_dep_data_22;
    assign token_22_34 = token_out_vec_22[16];

    // Process: write_back52_U0
    kernel_pr_hls_deadlock_detect_unit #(35, 23, 17, 17) kernel_pr_hls_deadlock_detect_unit_23 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_23),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_23),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_23),
        .token_in_vec(token_in_vec_23),
        .dl_detect_in(dl_detect_out),
        .origin(origin[23]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_23),
        .out_chan_dep_data(out_chan_dep_data_23),
        .token_out_vec(token_out_vec_23),
        .dl_detect_out(dl_in_vec[23]));

    assign proc_23_data_FIFO_blk[0] = 1'b0 | (~write_back52_U0.H_blk_n) | (~write_back52_U0.hyperedge_size_blk_n);
    assign proc_23_data_PIPO_blk[0] = 1'b0;
    assign proc_23_start_FIFO_blk[0] = 1'b0 | (~start_for_write_back52_U0_U.if_empty_n & write_back52_U0.ap_idle & ~start_for_write_back52_U0_U.if_write);
    assign proc_23_TLF_FIFO_blk[0] = 1'b0;
    assign proc_23_input_sync_blk[0] = 1'b0;
    assign proc_23_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_23[0] = dl_detect_out ? proc_dep_vld_vec_23_reg[0] : (proc_23_data_FIFO_blk[0] | proc_23_data_PIPO_blk[0] | proc_23_start_FIFO_blk[0] | proc_23_TLF_FIFO_blk[0] | proc_23_input_sync_blk[0] | proc_23_output_sync_blk[0]);
    assign proc_23_data_FIFO_blk[1] = 1'b0 | (~write_back52_U0.value_stream_V_V4_blk_n);
    assign proc_23_data_PIPO_blk[1] = 1'b0;
    assign proc_23_start_FIFO_blk[1] = 1'b0;
    assign proc_23_TLF_FIFO_blk[1] = 1'b0;
    assign proc_23_input_sync_blk[1] = 1'b0;
    assign proc_23_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_23[1] = dl_detect_out ? proc_dep_vld_vec_23_reg[1] : (proc_23_data_FIFO_blk[1] | proc_23_data_PIPO_blk[1] | proc_23_start_FIFO_blk[1] | proc_23_TLF_FIFO_blk[1] | proc_23_input_sync_blk[1] | proc_23_output_sync_blk[1]);
    assign proc_23_data_FIFO_blk[2] = 1'b0;
    assign proc_23_data_PIPO_blk[2] = 1'b0;
    assign proc_23_start_FIFO_blk[2] = 1'b0;
    assign proc_23_TLF_FIFO_blk[2] = 1'b0;
    assign proc_23_input_sync_blk[2] = 1'b0;
    assign proc_23_output_sync_blk[2] = 1'b0 | (ap_done_reg_4 & write_back52_U0.ap_done & ~write_back48_U0.ap_done);
    assign proc_dep_vld_vec_23[2] = dl_detect_out ? proc_dep_vld_vec_23_reg[2] : (proc_23_data_FIFO_blk[2] | proc_23_data_PIPO_blk[2] | proc_23_start_FIFO_blk[2] | proc_23_TLF_FIFO_blk[2] | proc_23_input_sync_blk[2] | proc_23_output_sync_blk[2]);
    assign proc_23_data_FIFO_blk[3] = 1'b0;
    assign proc_23_data_PIPO_blk[3] = 1'b0;
    assign proc_23_start_FIFO_blk[3] = 1'b0;
    assign proc_23_TLF_FIFO_blk[3] = 1'b0;
    assign proc_23_input_sync_blk[3] = 1'b0;
    assign proc_23_output_sync_blk[3] = 1'b0 | (ap_done_reg_4 & write_back52_U0.ap_done & ~write_back49_U0.ap_done);
    assign proc_dep_vld_vec_23[3] = dl_detect_out ? proc_dep_vld_vec_23_reg[3] : (proc_23_data_FIFO_blk[3] | proc_23_data_PIPO_blk[3] | proc_23_start_FIFO_blk[3] | proc_23_TLF_FIFO_blk[3] | proc_23_input_sync_blk[3] | proc_23_output_sync_blk[3]);
    assign proc_23_data_FIFO_blk[4] = 1'b0;
    assign proc_23_data_PIPO_blk[4] = 1'b0;
    assign proc_23_start_FIFO_blk[4] = 1'b0;
    assign proc_23_TLF_FIFO_blk[4] = 1'b0;
    assign proc_23_input_sync_blk[4] = 1'b0;
    assign proc_23_output_sync_blk[4] = 1'b0 | (ap_done_reg_4 & write_back52_U0.ap_done & ~write_back50_U0.ap_done);
    assign proc_dep_vld_vec_23[4] = dl_detect_out ? proc_dep_vld_vec_23_reg[4] : (proc_23_data_FIFO_blk[4] | proc_23_data_PIPO_blk[4] | proc_23_start_FIFO_blk[4] | proc_23_TLF_FIFO_blk[4] | proc_23_input_sync_blk[4] | proc_23_output_sync_blk[4]);
    assign proc_23_data_FIFO_blk[5] = 1'b0;
    assign proc_23_data_PIPO_blk[5] = 1'b0;
    assign proc_23_start_FIFO_blk[5] = 1'b0;
    assign proc_23_TLF_FIFO_blk[5] = 1'b0;
    assign proc_23_input_sync_blk[5] = 1'b0;
    assign proc_23_output_sync_blk[5] = 1'b0 | (ap_done_reg_4 & write_back52_U0.ap_done & ~write_back51_U0.ap_done);
    assign proc_dep_vld_vec_23[5] = dl_detect_out ? proc_dep_vld_vec_23_reg[5] : (proc_23_data_FIFO_blk[5] | proc_23_data_PIPO_blk[5] | proc_23_start_FIFO_blk[5] | proc_23_TLF_FIFO_blk[5] | proc_23_input_sync_blk[5] | proc_23_output_sync_blk[5]);
    assign proc_23_data_FIFO_blk[6] = 1'b0;
    assign proc_23_data_PIPO_blk[6] = 1'b0;
    assign proc_23_start_FIFO_blk[6] = 1'b0;
    assign proc_23_TLF_FIFO_blk[6] = 1'b0;
    assign proc_23_input_sync_blk[6] = 1'b0;
    assign proc_23_output_sync_blk[6] = 1'b0 | (ap_done_reg_4 & write_back52_U0.ap_done & ~write_back53_U0.ap_done);
    assign proc_dep_vld_vec_23[6] = dl_detect_out ? proc_dep_vld_vec_23_reg[6] : (proc_23_data_FIFO_blk[6] | proc_23_data_PIPO_blk[6] | proc_23_start_FIFO_blk[6] | proc_23_TLF_FIFO_blk[6] | proc_23_input_sync_blk[6] | proc_23_output_sync_blk[6]);
    assign proc_23_data_FIFO_blk[7] = 1'b0;
    assign proc_23_data_PIPO_blk[7] = 1'b0;
    assign proc_23_start_FIFO_blk[7] = 1'b0;
    assign proc_23_TLF_FIFO_blk[7] = 1'b0;
    assign proc_23_input_sync_blk[7] = 1'b0;
    assign proc_23_output_sync_blk[7] = 1'b0 | (ap_done_reg_4 & write_back52_U0.ap_done & ~write_back54_U0.ap_done);
    assign proc_dep_vld_vec_23[7] = dl_detect_out ? proc_dep_vld_vec_23_reg[7] : (proc_23_data_FIFO_blk[7] | proc_23_data_PIPO_blk[7] | proc_23_start_FIFO_blk[7] | proc_23_TLF_FIFO_blk[7] | proc_23_input_sync_blk[7] | proc_23_output_sync_blk[7]);
    assign proc_23_data_FIFO_blk[8] = 1'b0;
    assign proc_23_data_PIPO_blk[8] = 1'b0;
    assign proc_23_start_FIFO_blk[8] = 1'b0;
    assign proc_23_TLF_FIFO_blk[8] = 1'b0;
    assign proc_23_input_sync_blk[8] = 1'b0;
    assign proc_23_output_sync_blk[8] = 1'b0 | (ap_done_reg_4 & write_back52_U0.ap_done & ~write_back55_U0.ap_done);
    assign proc_dep_vld_vec_23[8] = dl_detect_out ? proc_dep_vld_vec_23_reg[8] : (proc_23_data_FIFO_blk[8] | proc_23_data_PIPO_blk[8] | proc_23_start_FIFO_blk[8] | proc_23_TLF_FIFO_blk[8] | proc_23_input_sync_blk[8] | proc_23_output_sync_blk[8]);
    assign proc_23_data_FIFO_blk[9] = 1'b0;
    assign proc_23_data_PIPO_blk[9] = 1'b0;
    assign proc_23_start_FIFO_blk[9] = 1'b0;
    assign proc_23_TLF_FIFO_blk[9] = 1'b0;
    assign proc_23_input_sync_blk[9] = 1'b0;
    assign proc_23_output_sync_blk[9] = 1'b0 | (ap_done_reg_4 & write_back52_U0.ap_done & ~write_back56_U0.ap_done);
    assign proc_dep_vld_vec_23[9] = dl_detect_out ? proc_dep_vld_vec_23_reg[9] : (proc_23_data_FIFO_blk[9] | proc_23_data_PIPO_blk[9] | proc_23_start_FIFO_blk[9] | proc_23_TLF_FIFO_blk[9] | proc_23_input_sync_blk[9] | proc_23_output_sync_blk[9]);
    assign proc_23_data_FIFO_blk[10] = 1'b0;
    assign proc_23_data_PIPO_blk[10] = 1'b0;
    assign proc_23_start_FIFO_blk[10] = 1'b0;
    assign proc_23_TLF_FIFO_blk[10] = 1'b0;
    assign proc_23_input_sync_blk[10] = 1'b0;
    assign proc_23_output_sync_blk[10] = 1'b0 | (ap_done_reg_4 & write_back52_U0.ap_done & ~write_back57_U0.ap_done);
    assign proc_dep_vld_vec_23[10] = dl_detect_out ? proc_dep_vld_vec_23_reg[10] : (proc_23_data_FIFO_blk[10] | proc_23_data_PIPO_blk[10] | proc_23_start_FIFO_blk[10] | proc_23_TLF_FIFO_blk[10] | proc_23_input_sync_blk[10] | proc_23_output_sync_blk[10]);
    assign proc_23_data_FIFO_blk[11] = 1'b0;
    assign proc_23_data_PIPO_blk[11] = 1'b0;
    assign proc_23_start_FIFO_blk[11] = 1'b0;
    assign proc_23_TLF_FIFO_blk[11] = 1'b0;
    assign proc_23_input_sync_blk[11] = 1'b0;
    assign proc_23_output_sync_blk[11] = 1'b0 | (ap_done_reg_4 & write_back52_U0.ap_done & ~write_back58_U0.ap_done);
    assign proc_dep_vld_vec_23[11] = dl_detect_out ? proc_dep_vld_vec_23_reg[11] : (proc_23_data_FIFO_blk[11] | proc_23_data_PIPO_blk[11] | proc_23_start_FIFO_blk[11] | proc_23_TLF_FIFO_blk[11] | proc_23_input_sync_blk[11] | proc_23_output_sync_blk[11]);
    assign proc_23_data_FIFO_blk[12] = 1'b0;
    assign proc_23_data_PIPO_blk[12] = 1'b0;
    assign proc_23_start_FIFO_blk[12] = 1'b0;
    assign proc_23_TLF_FIFO_blk[12] = 1'b0;
    assign proc_23_input_sync_blk[12] = 1'b0;
    assign proc_23_output_sync_blk[12] = 1'b0 | (ap_done_reg_4 & write_back52_U0.ap_done & ~write_back59_U0.ap_done);
    assign proc_dep_vld_vec_23[12] = dl_detect_out ? proc_dep_vld_vec_23_reg[12] : (proc_23_data_FIFO_blk[12] | proc_23_data_PIPO_blk[12] | proc_23_start_FIFO_blk[12] | proc_23_TLF_FIFO_blk[12] | proc_23_input_sync_blk[12] | proc_23_output_sync_blk[12]);
    assign proc_23_data_FIFO_blk[13] = 1'b0;
    assign proc_23_data_PIPO_blk[13] = 1'b0;
    assign proc_23_start_FIFO_blk[13] = 1'b0;
    assign proc_23_TLF_FIFO_blk[13] = 1'b0;
    assign proc_23_input_sync_blk[13] = 1'b0;
    assign proc_23_output_sync_blk[13] = 1'b0 | (ap_done_reg_4 & write_back52_U0.ap_done & ~write_back60_U0.ap_done);
    assign proc_dep_vld_vec_23[13] = dl_detect_out ? proc_dep_vld_vec_23_reg[13] : (proc_23_data_FIFO_blk[13] | proc_23_data_PIPO_blk[13] | proc_23_start_FIFO_blk[13] | proc_23_TLF_FIFO_blk[13] | proc_23_input_sync_blk[13] | proc_23_output_sync_blk[13]);
    assign proc_23_data_FIFO_blk[14] = 1'b0;
    assign proc_23_data_PIPO_blk[14] = 1'b0;
    assign proc_23_start_FIFO_blk[14] = 1'b0;
    assign proc_23_TLF_FIFO_blk[14] = 1'b0;
    assign proc_23_input_sync_blk[14] = 1'b0;
    assign proc_23_output_sync_blk[14] = 1'b0 | (ap_done_reg_4 & write_back52_U0.ap_done & ~write_back61_U0.ap_done);
    assign proc_dep_vld_vec_23[14] = dl_detect_out ? proc_dep_vld_vec_23_reg[14] : (proc_23_data_FIFO_blk[14] | proc_23_data_PIPO_blk[14] | proc_23_start_FIFO_blk[14] | proc_23_TLF_FIFO_blk[14] | proc_23_input_sync_blk[14] | proc_23_output_sync_blk[14]);
    assign proc_23_data_FIFO_blk[15] = 1'b0;
    assign proc_23_data_PIPO_blk[15] = 1'b0;
    assign proc_23_start_FIFO_blk[15] = 1'b0;
    assign proc_23_TLF_FIFO_blk[15] = 1'b0;
    assign proc_23_input_sync_blk[15] = 1'b0;
    assign proc_23_output_sync_blk[15] = 1'b0 | (ap_done_reg_4 & write_back52_U0.ap_done & ~write_back62_U0.ap_done);
    assign proc_dep_vld_vec_23[15] = dl_detect_out ? proc_dep_vld_vec_23_reg[15] : (proc_23_data_FIFO_blk[15] | proc_23_data_PIPO_blk[15] | proc_23_start_FIFO_blk[15] | proc_23_TLF_FIFO_blk[15] | proc_23_input_sync_blk[15] | proc_23_output_sync_blk[15]);
    assign proc_23_data_FIFO_blk[16] = 1'b0;
    assign proc_23_data_PIPO_blk[16] = 1'b0;
    assign proc_23_start_FIFO_blk[16] = 1'b0;
    assign proc_23_TLF_FIFO_blk[16] = 1'b0;
    assign proc_23_input_sync_blk[16] = 1'b0;
    assign proc_23_output_sync_blk[16] = 1'b0 | (ap_done_reg_4 & write_back52_U0.ap_done & ~write_back63_U0.ap_done);
    assign proc_dep_vld_vec_23[16] = dl_detect_out ? proc_dep_vld_vec_23_reg[16] : (proc_23_data_FIFO_blk[16] | proc_23_data_PIPO_blk[16] | proc_23_start_FIFO_blk[16] | proc_23_TLF_FIFO_blk[16] | proc_23_input_sync_blk[16] | proc_23_output_sync_blk[16]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_23_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_23_reg <= proc_dep_vld_vec_23;
        end
    end
    assign in_chan_dep_vld_vec_23[0] = dep_chan_vld_0_23;
    assign in_chan_dep_data_vec_23[34 : 0] = dep_chan_data_0_23;
    assign token_in_vec_23[0] = token_0_23;
    assign in_chan_dep_vld_vec_23[1] = dep_chan_vld_7_23;
    assign in_chan_dep_data_vec_23[69 : 35] = dep_chan_data_7_23;
    assign token_in_vec_23[1] = token_7_23;
    assign in_chan_dep_vld_vec_23[2] = dep_chan_vld_19_23;
    assign in_chan_dep_data_vec_23[104 : 70] = dep_chan_data_19_23;
    assign token_in_vec_23[2] = token_19_23;
    assign in_chan_dep_vld_vec_23[3] = dep_chan_vld_20_23;
    assign in_chan_dep_data_vec_23[139 : 105] = dep_chan_data_20_23;
    assign token_in_vec_23[3] = token_20_23;
    assign in_chan_dep_vld_vec_23[4] = dep_chan_vld_21_23;
    assign in_chan_dep_data_vec_23[174 : 140] = dep_chan_data_21_23;
    assign token_in_vec_23[4] = token_21_23;
    assign in_chan_dep_vld_vec_23[5] = dep_chan_vld_22_23;
    assign in_chan_dep_data_vec_23[209 : 175] = dep_chan_data_22_23;
    assign token_in_vec_23[5] = token_22_23;
    assign in_chan_dep_vld_vec_23[6] = dep_chan_vld_24_23;
    assign in_chan_dep_data_vec_23[244 : 210] = dep_chan_data_24_23;
    assign token_in_vec_23[6] = token_24_23;
    assign in_chan_dep_vld_vec_23[7] = dep_chan_vld_25_23;
    assign in_chan_dep_data_vec_23[279 : 245] = dep_chan_data_25_23;
    assign token_in_vec_23[7] = token_25_23;
    assign in_chan_dep_vld_vec_23[8] = dep_chan_vld_26_23;
    assign in_chan_dep_data_vec_23[314 : 280] = dep_chan_data_26_23;
    assign token_in_vec_23[8] = token_26_23;
    assign in_chan_dep_vld_vec_23[9] = dep_chan_vld_27_23;
    assign in_chan_dep_data_vec_23[349 : 315] = dep_chan_data_27_23;
    assign token_in_vec_23[9] = token_27_23;
    assign in_chan_dep_vld_vec_23[10] = dep_chan_vld_28_23;
    assign in_chan_dep_data_vec_23[384 : 350] = dep_chan_data_28_23;
    assign token_in_vec_23[10] = token_28_23;
    assign in_chan_dep_vld_vec_23[11] = dep_chan_vld_29_23;
    assign in_chan_dep_data_vec_23[419 : 385] = dep_chan_data_29_23;
    assign token_in_vec_23[11] = token_29_23;
    assign in_chan_dep_vld_vec_23[12] = dep_chan_vld_30_23;
    assign in_chan_dep_data_vec_23[454 : 420] = dep_chan_data_30_23;
    assign token_in_vec_23[12] = token_30_23;
    assign in_chan_dep_vld_vec_23[13] = dep_chan_vld_31_23;
    assign in_chan_dep_data_vec_23[489 : 455] = dep_chan_data_31_23;
    assign token_in_vec_23[13] = token_31_23;
    assign in_chan_dep_vld_vec_23[14] = dep_chan_vld_32_23;
    assign in_chan_dep_data_vec_23[524 : 490] = dep_chan_data_32_23;
    assign token_in_vec_23[14] = token_32_23;
    assign in_chan_dep_vld_vec_23[15] = dep_chan_vld_33_23;
    assign in_chan_dep_data_vec_23[559 : 525] = dep_chan_data_33_23;
    assign token_in_vec_23[15] = token_33_23;
    assign in_chan_dep_vld_vec_23[16] = dep_chan_vld_34_23;
    assign in_chan_dep_data_vec_23[594 : 560] = dep_chan_data_34_23;
    assign token_in_vec_23[16] = token_34_23;
    assign dep_chan_vld_23_0 = out_chan_dep_vld_vec_23[0];
    assign dep_chan_data_23_0 = out_chan_dep_data_23;
    assign token_23_0 = token_out_vec_23[0];
    assign dep_chan_vld_23_7 = out_chan_dep_vld_vec_23[1];
    assign dep_chan_data_23_7 = out_chan_dep_data_23;
    assign token_23_7 = token_out_vec_23[1];
    assign dep_chan_vld_23_19 = out_chan_dep_vld_vec_23[2];
    assign dep_chan_data_23_19 = out_chan_dep_data_23;
    assign token_23_19 = token_out_vec_23[2];
    assign dep_chan_vld_23_20 = out_chan_dep_vld_vec_23[3];
    assign dep_chan_data_23_20 = out_chan_dep_data_23;
    assign token_23_20 = token_out_vec_23[3];
    assign dep_chan_vld_23_21 = out_chan_dep_vld_vec_23[4];
    assign dep_chan_data_23_21 = out_chan_dep_data_23;
    assign token_23_21 = token_out_vec_23[4];
    assign dep_chan_vld_23_22 = out_chan_dep_vld_vec_23[5];
    assign dep_chan_data_23_22 = out_chan_dep_data_23;
    assign token_23_22 = token_out_vec_23[5];
    assign dep_chan_vld_23_24 = out_chan_dep_vld_vec_23[6];
    assign dep_chan_data_23_24 = out_chan_dep_data_23;
    assign token_23_24 = token_out_vec_23[6];
    assign dep_chan_vld_23_25 = out_chan_dep_vld_vec_23[7];
    assign dep_chan_data_23_25 = out_chan_dep_data_23;
    assign token_23_25 = token_out_vec_23[7];
    assign dep_chan_vld_23_26 = out_chan_dep_vld_vec_23[8];
    assign dep_chan_data_23_26 = out_chan_dep_data_23;
    assign token_23_26 = token_out_vec_23[8];
    assign dep_chan_vld_23_27 = out_chan_dep_vld_vec_23[9];
    assign dep_chan_data_23_27 = out_chan_dep_data_23;
    assign token_23_27 = token_out_vec_23[9];
    assign dep_chan_vld_23_28 = out_chan_dep_vld_vec_23[10];
    assign dep_chan_data_23_28 = out_chan_dep_data_23;
    assign token_23_28 = token_out_vec_23[10];
    assign dep_chan_vld_23_29 = out_chan_dep_vld_vec_23[11];
    assign dep_chan_data_23_29 = out_chan_dep_data_23;
    assign token_23_29 = token_out_vec_23[11];
    assign dep_chan_vld_23_30 = out_chan_dep_vld_vec_23[12];
    assign dep_chan_data_23_30 = out_chan_dep_data_23;
    assign token_23_30 = token_out_vec_23[12];
    assign dep_chan_vld_23_31 = out_chan_dep_vld_vec_23[13];
    assign dep_chan_data_23_31 = out_chan_dep_data_23;
    assign token_23_31 = token_out_vec_23[13];
    assign dep_chan_vld_23_32 = out_chan_dep_vld_vec_23[14];
    assign dep_chan_data_23_32 = out_chan_dep_data_23;
    assign token_23_32 = token_out_vec_23[14];
    assign dep_chan_vld_23_33 = out_chan_dep_vld_vec_23[15];
    assign dep_chan_data_23_33 = out_chan_dep_data_23;
    assign token_23_33 = token_out_vec_23[15];
    assign dep_chan_vld_23_34 = out_chan_dep_vld_vec_23[16];
    assign dep_chan_data_23_34 = out_chan_dep_data_23;
    assign token_23_34 = token_out_vec_23[16];

    // Process: write_back53_U0
    kernel_pr_hls_deadlock_detect_unit #(35, 24, 17, 17) kernel_pr_hls_deadlock_detect_unit_24 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_24),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_24),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_24),
        .token_in_vec(token_in_vec_24),
        .dl_detect_in(dl_detect_out),
        .origin(origin[24]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_24),
        .out_chan_dep_data(out_chan_dep_data_24),
        .token_out_vec(token_out_vec_24),
        .dl_detect_out(dl_in_vec[24]));

    assign proc_24_data_FIFO_blk[0] = 1'b0 | (~write_back53_U0.H_blk_n) | (~write_back53_U0.hyperedge_size_blk_n);
    assign proc_24_data_PIPO_blk[0] = 1'b0;
    assign proc_24_start_FIFO_blk[0] = 1'b0 | (~start_for_write_back53_U0_U.if_empty_n & write_back53_U0.ap_idle & ~start_for_write_back53_U0_U.if_write);
    assign proc_24_TLF_FIFO_blk[0] = 1'b0;
    assign proc_24_input_sync_blk[0] = 1'b0;
    assign proc_24_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_24[0] = dl_detect_out ? proc_dep_vld_vec_24_reg[0] : (proc_24_data_FIFO_blk[0] | proc_24_data_PIPO_blk[0] | proc_24_start_FIFO_blk[0] | proc_24_TLF_FIFO_blk[0] | proc_24_input_sync_blk[0] | proc_24_output_sync_blk[0]);
    assign proc_24_data_FIFO_blk[1] = 1'b0 | (~write_back53_U0.value_stream_V_V5_blk_n);
    assign proc_24_data_PIPO_blk[1] = 1'b0;
    assign proc_24_start_FIFO_blk[1] = 1'b0;
    assign proc_24_TLF_FIFO_blk[1] = 1'b0;
    assign proc_24_input_sync_blk[1] = 1'b0;
    assign proc_24_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_24[1] = dl_detect_out ? proc_dep_vld_vec_24_reg[1] : (proc_24_data_FIFO_blk[1] | proc_24_data_PIPO_blk[1] | proc_24_start_FIFO_blk[1] | proc_24_TLF_FIFO_blk[1] | proc_24_input_sync_blk[1] | proc_24_output_sync_blk[1]);
    assign proc_24_data_FIFO_blk[2] = 1'b0;
    assign proc_24_data_PIPO_blk[2] = 1'b0;
    assign proc_24_start_FIFO_blk[2] = 1'b0;
    assign proc_24_TLF_FIFO_blk[2] = 1'b0;
    assign proc_24_input_sync_blk[2] = 1'b0;
    assign proc_24_output_sync_blk[2] = 1'b0 | (ap_done_reg_5 & write_back53_U0.ap_done & ~write_back48_U0.ap_done);
    assign proc_dep_vld_vec_24[2] = dl_detect_out ? proc_dep_vld_vec_24_reg[2] : (proc_24_data_FIFO_blk[2] | proc_24_data_PIPO_blk[2] | proc_24_start_FIFO_blk[2] | proc_24_TLF_FIFO_blk[2] | proc_24_input_sync_blk[2] | proc_24_output_sync_blk[2]);
    assign proc_24_data_FIFO_blk[3] = 1'b0;
    assign proc_24_data_PIPO_blk[3] = 1'b0;
    assign proc_24_start_FIFO_blk[3] = 1'b0;
    assign proc_24_TLF_FIFO_blk[3] = 1'b0;
    assign proc_24_input_sync_blk[3] = 1'b0;
    assign proc_24_output_sync_blk[3] = 1'b0 | (ap_done_reg_5 & write_back53_U0.ap_done & ~write_back49_U0.ap_done);
    assign proc_dep_vld_vec_24[3] = dl_detect_out ? proc_dep_vld_vec_24_reg[3] : (proc_24_data_FIFO_blk[3] | proc_24_data_PIPO_blk[3] | proc_24_start_FIFO_blk[3] | proc_24_TLF_FIFO_blk[3] | proc_24_input_sync_blk[3] | proc_24_output_sync_blk[3]);
    assign proc_24_data_FIFO_blk[4] = 1'b0;
    assign proc_24_data_PIPO_blk[4] = 1'b0;
    assign proc_24_start_FIFO_blk[4] = 1'b0;
    assign proc_24_TLF_FIFO_blk[4] = 1'b0;
    assign proc_24_input_sync_blk[4] = 1'b0;
    assign proc_24_output_sync_blk[4] = 1'b0 | (ap_done_reg_5 & write_back53_U0.ap_done & ~write_back50_U0.ap_done);
    assign proc_dep_vld_vec_24[4] = dl_detect_out ? proc_dep_vld_vec_24_reg[4] : (proc_24_data_FIFO_blk[4] | proc_24_data_PIPO_blk[4] | proc_24_start_FIFO_blk[4] | proc_24_TLF_FIFO_blk[4] | proc_24_input_sync_blk[4] | proc_24_output_sync_blk[4]);
    assign proc_24_data_FIFO_blk[5] = 1'b0;
    assign proc_24_data_PIPO_blk[5] = 1'b0;
    assign proc_24_start_FIFO_blk[5] = 1'b0;
    assign proc_24_TLF_FIFO_blk[5] = 1'b0;
    assign proc_24_input_sync_blk[5] = 1'b0;
    assign proc_24_output_sync_blk[5] = 1'b0 | (ap_done_reg_5 & write_back53_U0.ap_done & ~write_back51_U0.ap_done);
    assign proc_dep_vld_vec_24[5] = dl_detect_out ? proc_dep_vld_vec_24_reg[5] : (proc_24_data_FIFO_blk[5] | proc_24_data_PIPO_blk[5] | proc_24_start_FIFO_blk[5] | proc_24_TLF_FIFO_blk[5] | proc_24_input_sync_blk[5] | proc_24_output_sync_blk[5]);
    assign proc_24_data_FIFO_blk[6] = 1'b0;
    assign proc_24_data_PIPO_blk[6] = 1'b0;
    assign proc_24_start_FIFO_blk[6] = 1'b0;
    assign proc_24_TLF_FIFO_blk[6] = 1'b0;
    assign proc_24_input_sync_blk[6] = 1'b0;
    assign proc_24_output_sync_blk[6] = 1'b0 | (ap_done_reg_5 & write_back53_U0.ap_done & ~write_back52_U0.ap_done);
    assign proc_dep_vld_vec_24[6] = dl_detect_out ? proc_dep_vld_vec_24_reg[6] : (proc_24_data_FIFO_blk[6] | proc_24_data_PIPO_blk[6] | proc_24_start_FIFO_blk[6] | proc_24_TLF_FIFO_blk[6] | proc_24_input_sync_blk[6] | proc_24_output_sync_blk[6]);
    assign proc_24_data_FIFO_blk[7] = 1'b0;
    assign proc_24_data_PIPO_blk[7] = 1'b0;
    assign proc_24_start_FIFO_blk[7] = 1'b0;
    assign proc_24_TLF_FIFO_blk[7] = 1'b0;
    assign proc_24_input_sync_blk[7] = 1'b0;
    assign proc_24_output_sync_blk[7] = 1'b0 | (ap_done_reg_5 & write_back53_U0.ap_done & ~write_back54_U0.ap_done);
    assign proc_dep_vld_vec_24[7] = dl_detect_out ? proc_dep_vld_vec_24_reg[7] : (proc_24_data_FIFO_blk[7] | proc_24_data_PIPO_blk[7] | proc_24_start_FIFO_blk[7] | proc_24_TLF_FIFO_blk[7] | proc_24_input_sync_blk[7] | proc_24_output_sync_blk[7]);
    assign proc_24_data_FIFO_blk[8] = 1'b0;
    assign proc_24_data_PIPO_blk[8] = 1'b0;
    assign proc_24_start_FIFO_blk[8] = 1'b0;
    assign proc_24_TLF_FIFO_blk[8] = 1'b0;
    assign proc_24_input_sync_blk[8] = 1'b0;
    assign proc_24_output_sync_blk[8] = 1'b0 | (ap_done_reg_5 & write_back53_U0.ap_done & ~write_back55_U0.ap_done);
    assign proc_dep_vld_vec_24[8] = dl_detect_out ? proc_dep_vld_vec_24_reg[8] : (proc_24_data_FIFO_blk[8] | proc_24_data_PIPO_blk[8] | proc_24_start_FIFO_blk[8] | proc_24_TLF_FIFO_blk[8] | proc_24_input_sync_blk[8] | proc_24_output_sync_blk[8]);
    assign proc_24_data_FIFO_blk[9] = 1'b0;
    assign proc_24_data_PIPO_blk[9] = 1'b0;
    assign proc_24_start_FIFO_blk[9] = 1'b0;
    assign proc_24_TLF_FIFO_blk[9] = 1'b0;
    assign proc_24_input_sync_blk[9] = 1'b0;
    assign proc_24_output_sync_blk[9] = 1'b0 | (ap_done_reg_5 & write_back53_U0.ap_done & ~write_back56_U0.ap_done);
    assign proc_dep_vld_vec_24[9] = dl_detect_out ? proc_dep_vld_vec_24_reg[9] : (proc_24_data_FIFO_blk[9] | proc_24_data_PIPO_blk[9] | proc_24_start_FIFO_blk[9] | proc_24_TLF_FIFO_blk[9] | proc_24_input_sync_blk[9] | proc_24_output_sync_blk[9]);
    assign proc_24_data_FIFO_blk[10] = 1'b0;
    assign proc_24_data_PIPO_blk[10] = 1'b0;
    assign proc_24_start_FIFO_blk[10] = 1'b0;
    assign proc_24_TLF_FIFO_blk[10] = 1'b0;
    assign proc_24_input_sync_blk[10] = 1'b0;
    assign proc_24_output_sync_blk[10] = 1'b0 | (ap_done_reg_5 & write_back53_U0.ap_done & ~write_back57_U0.ap_done);
    assign proc_dep_vld_vec_24[10] = dl_detect_out ? proc_dep_vld_vec_24_reg[10] : (proc_24_data_FIFO_blk[10] | proc_24_data_PIPO_blk[10] | proc_24_start_FIFO_blk[10] | proc_24_TLF_FIFO_blk[10] | proc_24_input_sync_blk[10] | proc_24_output_sync_blk[10]);
    assign proc_24_data_FIFO_blk[11] = 1'b0;
    assign proc_24_data_PIPO_blk[11] = 1'b0;
    assign proc_24_start_FIFO_blk[11] = 1'b0;
    assign proc_24_TLF_FIFO_blk[11] = 1'b0;
    assign proc_24_input_sync_blk[11] = 1'b0;
    assign proc_24_output_sync_blk[11] = 1'b0 | (ap_done_reg_5 & write_back53_U0.ap_done & ~write_back58_U0.ap_done);
    assign proc_dep_vld_vec_24[11] = dl_detect_out ? proc_dep_vld_vec_24_reg[11] : (proc_24_data_FIFO_blk[11] | proc_24_data_PIPO_blk[11] | proc_24_start_FIFO_blk[11] | proc_24_TLF_FIFO_blk[11] | proc_24_input_sync_blk[11] | proc_24_output_sync_blk[11]);
    assign proc_24_data_FIFO_blk[12] = 1'b0;
    assign proc_24_data_PIPO_blk[12] = 1'b0;
    assign proc_24_start_FIFO_blk[12] = 1'b0;
    assign proc_24_TLF_FIFO_blk[12] = 1'b0;
    assign proc_24_input_sync_blk[12] = 1'b0;
    assign proc_24_output_sync_blk[12] = 1'b0 | (ap_done_reg_5 & write_back53_U0.ap_done & ~write_back59_U0.ap_done);
    assign proc_dep_vld_vec_24[12] = dl_detect_out ? proc_dep_vld_vec_24_reg[12] : (proc_24_data_FIFO_blk[12] | proc_24_data_PIPO_blk[12] | proc_24_start_FIFO_blk[12] | proc_24_TLF_FIFO_blk[12] | proc_24_input_sync_blk[12] | proc_24_output_sync_blk[12]);
    assign proc_24_data_FIFO_blk[13] = 1'b0;
    assign proc_24_data_PIPO_blk[13] = 1'b0;
    assign proc_24_start_FIFO_blk[13] = 1'b0;
    assign proc_24_TLF_FIFO_blk[13] = 1'b0;
    assign proc_24_input_sync_blk[13] = 1'b0;
    assign proc_24_output_sync_blk[13] = 1'b0 | (ap_done_reg_5 & write_back53_U0.ap_done & ~write_back60_U0.ap_done);
    assign proc_dep_vld_vec_24[13] = dl_detect_out ? proc_dep_vld_vec_24_reg[13] : (proc_24_data_FIFO_blk[13] | proc_24_data_PIPO_blk[13] | proc_24_start_FIFO_blk[13] | proc_24_TLF_FIFO_blk[13] | proc_24_input_sync_blk[13] | proc_24_output_sync_blk[13]);
    assign proc_24_data_FIFO_blk[14] = 1'b0;
    assign proc_24_data_PIPO_blk[14] = 1'b0;
    assign proc_24_start_FIFO_blk[14] = 1'b0;
    assign proc_24_TLF_FIFO_blk[14] = 1'b0;
    assign proc_24_input_sync_blk[14] = 1'b0;
    assign proc_24_output_sync_blk[14] = 1'b0 | (ap_done_reg_5 & write_back53_U0.ap_done & ~write_back61_U0.ap_done);
    assign proc_dep_vld_vec_24[14] = dl_detect_out ? proc_dep_vld_vec_24_reg[14] : (proc_24_data_FIFO_blk[14] | proc_24_data_PIPO_blk[14] | proc_24_start_FIFO_blk[14] | proc_24_TLF_FIFO_blk[14] | proc_24_input_sync_blk[14] | proc_24_output_sync_blk[14]);
    assign proc_24_data_FIFO_blk[15] = 1'b0;
    assign proc_24_data_PIPO_blk[15] = 1'b0;
    assign proc_24_start_FIFO_blk[15] = 1'b0;
    assign proc_24_TLF_FIFO_blk[15] = 1'b0;
    assign proc_24_input_sync_blk[15] = 1'b0;
    assign proc_24_output_sync_blk[15] = 1'b0 | (ap_done_reg_5 & write_back53_U0.ap_done & ~write_back62_U0.ap_done);
    assign proc_dep_vld_vec_24[15] = dl_detect_out ? proc_dep_vld_vec_24_reg[15] : (proc_24_data_FIFO_blk[15] | proc_24_data_PIPO_blk[15] | proc_24_start_FIFO_blk[15] | proc_24_TLF_FIFO_blk[15] | proc_24_input_sync_blk[15] | proc_24_output_sync_blk[15]);
    assign proc_24_data_FIFO_blk[16] = 1'b0;
    assign proc_24_data_PIPO_blk[16] = 1'b0;
    assign proc_24_start_FIFO_blk[16] = 1'b0;
    assign proc_24_TLF_FIFO_blk[16] = 1'b0;
    assign proc_24_input_sync_blk[16] = 1'b0;
    assign proc_24_output_sync_blk[16] = 1'b0 | (ap_done_reg_5 & write_back53_U0.ap_done & ~write_back63_U0.ap_done);
    assign proc_dep_vld_vec_24[16] = dl_detect_out ? proc_dep_vld_vec_24_reg[16] : (proc_24_data_FIFO_blk[16] | proc_24_data_PIPO_blk[16] | proc_24_start_FIFO_blk[16] | proc_24_TLF_FIFO_blk[16] | proc_24_input_sync_blk[16] | proc_24_output_sync_blk[16]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_24_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_24_reg <= proc_dep_vld_vec_24;
        end
    end
    assign in_chan_dep_vld_vec_24[0] = dep_chan_vld_0_24;
    assign in_chan_dep_data_vec_24[34 : 0] = dep_chan_data_0_24;
    assign token_in_vec_24[0] = token_0_24;
    assign in_chan_dep_vld_vec_24[1] = dep_chan_vld_8_24;
    assign in_chan_dep_data_vec_24[69 : 35] = dep_chan_data_8_24;
    assign token_in_vec_24[1] = token_8_24;
    assign in_chan_dep_vld_vec_24[2] = dep_chan_vld_19_24;
    assign in_chan_dep_data_vec_24[104 : 70] = dep_chan_data_19_24;
    assign token_in_vec_24[2] = token_19_24;
    assign in_chan_dep_vld_vec_24[3] = dep_chan_vld_20_24;
    assign in_chan_dep_data_vec_24[139 : 105] = dep_chan_data_20_24;
    assign token_in_vec_24[3] = token_20_24;
    assign in_chan_dep_vld_vec_24[4] = dep_chan_vld_21_24;
    assign in_chan_dep_data_vec_24[174 : 140] = dep_chan_data_21_24;
    assign token_in_vec_24[4] = token_21_24;
    assign in_chan_dep_vld_vec_24[5] = dep_chan_vld_22_24;
    assign in_chan_dep_data_vec_24[209 : 175] = dep_chan_data_22_24;
    assign token_in_vec_24[5] = token_22_24;
    assign in_chan_dep_vld_vec_24[6] = dep_chan_vld_23_24;
    assign in_chan_dep_data_vec_24[244 : 210] = dep_chan_data_23_24;
    assign token_in_vec_24[6] = token_23_24;
    assign in_chan_dep_vld_vec_24[7] = dep_chan_vld_25_24;
    assign in_chan_dep_data_vec_24[279 : 245] = dep_chan_data_25_24;
    assign token_in_vec_24[7] = token_25_24;
    assign in_chan_dep_vld_vec_24[8] = dep_chan_vld_26_24;
    assign in_chan_dep_data_vec_24[314 : 280] = dep_chan_data_26_24;
    assign token_in_vec_24[8] = token_26_24;
    assign in_chan_dep_vld_vec_24[9] = dep_chan_vld_27_24;
    assign in_chan_dep_data_vec_24[349 : 315] = dep_chan_data_27_24;
    assign token_in_vec_24[9] = token_27_24;
    assign in_chan_dep_vld_vec_24[10] = dep_chan_vld_28_24;
    assign in_chan_dep_data_vec_24[384 : 350] = dep_chan_data_28_24;
    assign token_in_vec_24[10] = token_28_24;
    assign in_chan_dep_vld_vec_24[11] = dep_chan_vld_29_24;
    assign in_chan_dep_data_vec_24[419 : 385] = dep_chan_data_29_24;
    assign token_in_vec_24[11] = token_29_24;
    assign in_chan_dep_vld_vec_24[12] = dep_chan_vld_30_24;
    assign in_chan_dep_data_vec_24[454 : 420] = dep_chan_data_30_24;
    assign token_in_vec_24[12] = token_30_24;
    assign in_chan_dep_vld_vec_24[13] = dep_chan_vld_31_24;
    assign in_chan_dep_data_vec_24[489 : 455] = dep_chan_data_31_24;
    assign token_in_vec_24[13] = token_31_24;
    assign in_chan_dep_vld_vec_24[14] = dep_chan_vld_32_24;
    assign in_chan_dep_data_vec_24[524 : 490] = dep_chan_data_32_24;
    assign token_in_vec_24[14] = token_32_24;
    assign in_chan_dep_vld_vec_24[15] = dep_chan_vld_33_24;
    assign in_chan_dep_data_vec_24[559 : 525] = dep_chan_data_33_24;
    assign token_in_vec_24[15] = token_33_24;
    assign in_chan_dep_vld_vec_24[16] = dep_chan_vld_34_24;
    assign in_chan_dep_data_vec_24[594 : 560] = dep_chan_data_34_24;
    assign token_in_vec_24[16] = token_34_24;
    assign dep_chan_vld_24_0 = out_chan_dep_vld_vec_24[0];
    assign dep_chan_data_24_0 = out_chan_dep_data_24;
    assign token_24_0 = token_out_vec_24[0];
    assign dep_chan_vld_24_8 = out_chan_dep_vld_vec_24[1];
    assign dep_chan_data_24_8 = out_chan_dep_data_24;
    assign token_24_8 = token_out_vec_24[1];
    assign dep_chan_vld_24_19 = out_chan_dep_vld_vec_24[2];
    assign dep_chan_data_24_19 = out_chan_dep_data_24;
    assign token_24_19 = token_out_vec_24[2];
    assign dep_chan_vld_24_20 = out_chan_dep_vld_vec_24[3];
    assign dep_chan_data_24_20 = out_chan_dep_data_24;
    assign token_24_20 = token_out_vec_24[3];
    assign dep_chan_vld_24_21 = out_chan_dep_vld_vec_24[4];
    assign dep_chan_data_24_21 = out_chan_dep_data_24;
    assign token_24_21 = token_out_vec_24[4];
    assign dep_chan_vld_24_22 = out_chan_dep_vld_vec_24[5];
    assign dep_chan_data_24_22 = out_chan_dep_data_24;
    assign token_24_22 = token_out_vec_24[5];
    assign dep_chan_vld_24_23 = out_chan_dep_vld_vec_24[6];
    assign dep_chan_data_24_23 = out_chan_dep_data_24;
    assign token_24_23 = token_out_vec_24[6];
    assign dep_chan_vld_24_25 = out_chan_dep_vld_vec_24[7];
    assign dep_chan_data_24_25 = out_chan_dep_data_24;
    assign token_24_25 = token_out_vec_24[7];
    assign dep_chan_vld_24_26 = out_chan_dep_vld_vec_24[8];
    assign dep_chan_data_24_26 = out_chan_dep_data_24;
    assign token_24_26 = token_out_vec_24[8];
    assign dep_chan_vld_24_27 = out_chan_dep_vld_vec_24[9];
    assign dep_chan_data_24_27 = out_chan_dep_data_24;
    assign token_24_27 = token_out_vec_24[9];
    assign dep_chan_vld_24_28 = out_chan_dep_vld_vec_24[10];
    assign dep_chan_data_24_28 = out_chan_dep_data_24;
    assign token_24_28 = token_out_vec_24[10];
    assign dep_chan_vld_24_29 = out_chan_dep_vld_vec_24[11];
    assign dep_chan_data_24_29 = out_chan_dep_data_24;
    assign token_24_29 = token_out_vec_24[11];
    assign dep_chan_vld_24_30 = out_chan_dep_vld_vec_24[12];
    assign dep_chan_data_24_30 = out_chan_dep_data_24;
    assign token_24_30 = token_out_vec_24[12];
    assign dep_chan_vld_24_31 = out_chan_dep_vld_vec_24[13];
    assign dep_chan_data_24_31 = out_chan_dep_data_24;
    assign token_24_31 = token_out_vec_24[13];
    assign dep_chan_vld_24_32 = out_chan_dep_vld_vec_24[14];
    assign dep_chan_data_24_32 = out_chan_dep_data_24;
    assign token_24_32 = token_out_vec_24[14];
    assign dep_chan_vld_24_33 = out_chan_dep_vld_vec_24[15];
    assign dep_chan_data_24_33 = out_chan_dep_data_24;
    assign token_24_33 = token_out_vec_24[15];
    assign dep_chan_vld_24_34 = out_chan_dep_vld_vec_24[16];
    assign dep_chan_data_24_34 = out_chan_dep_data_24;
    assign token_24_34 = token_out_vec_24[16];

    // Process: write_back54_U0
    kernel_pr_hls_deadlock_detect_unit #(35, 25, 17, 17) kernel_pr_hls_deadlock_detect_unit_25 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_25),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_25),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_25),
        .token_in_vec(token_in_vec_25),
        .dl_detect_in(dl_detect_out),
        .origin(origin[25]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_25),
        .out_chan_dep_data(out_chan_dep_data_25),
        .token_out_vec(token_out_vec_25),
        .dl_detect_out(dl_in_vec[25]));

    assign proc_25_data_FIFO_blk[0] = 1'b0 | (~write_back54_U0.H_blk_n) | (~write_back54_U0.hyperedge_size_blk_n);
    assign proc_25_data_PIPO_blk[0] = 1'b0;
    assign proc_25_start_FIFO_blk[0] = 1'b0 | (~start_for_write_back54_U0_U.if_empty_n & write_back54_U0.ap_idle & ~start_for_write_back54_U0_U.if_write);
    assign proc_25_TLF_FIFO_blk[0] = 1'b0;
    assign proc_25_input_sync_blk[0] = 1'b0;
    assign proc_25_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_25[0] = dl_detect_out ? proc_dep_vld_vec_25_reg[0] : (proc_25_data_FIFO_blk[0] | proc_25_data_PIPO_blk[0] | proc_25_start_FIFO_blk[0] | proc_25_TLF_FIFO_blk[0] | proc_25_input_sync_blk[0] | proc_25_output_sync_blk[0]);
    assign proc_25_data_FIFO_blk[1] = 1'b0 | (~write_back54_U0.value_stream_V_V6_blk_n);
    assign proc_25_data_PIPO_blk[1] = 1'b0;
    assign proc_25_start_FIFO_blk[1] = 1'b0;
    assign proc_25_TLF_FIFO_blk[1] = 1'b0;
    assign proc_25_input_sync_blk[1] = 1'b0;
    assign proc_25_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_25[1] = dl_detect_out ? proc_dep_vld_vec_25_reg[1] : (proc_25_data_FIFO_blk[1] | proc_25_data_PIPO_blk[1] | proc_25_start_FIFO_blk[1] | proc_25_TLF_FIFO_blk[1] | proc_25_input_sync_blk[1] | proc_25_output_sync_blk[1]);
    assign proc_25_data_FIFO_blk[2] = 1'b0;
    assign proc_25_data_PIPO_blk[2] = 1'b0;
    assign proc_25_start_FIFO_blk[2] = 1'b0;
    assign proc_25_TLF_FIFO_blk[2] = 1'b0;
    assign proc_25_input_sync_blk[2] = 1'b0;
    assign proc_25_output_sync_blk[2] = 1'b0 | (ap_done_reg_6 & write_back54_U0.ap_done & ~write_back48_U0.ap_done);
    assign proc_dep_vld_vec_25[2] = dl_detect_out ? proc_dep_vld_vec_25_reg[2] : (proc_25_data_FIFO_blk[2] | proc_25_data_PIPO_blk[2] | proc_25_start_FIFO_blk[2] | proc_25_TLF_FIFO_blk[2] | proc_25_input_sync_blk[2] | proc_25_output_sync_blk[2]);
    assign proc_25_data_FIFO_blk[3] = 1'b0;
    assign proc_25_data_PIPO_blk[3] = 1'b0;
    assign proc_25_start_FIFO_blk[3] = 1'b0;
    assign proc_25_TLF_FIFO_blk[3] = 1'b0;
    assign proc_25_input_sync_blk[3] = 1'b0;
    assign proc_25_output_sync_blk[3] = 1'b0 | (ap_done_reg_6 & write_back54_U0.ap_done & ~write_back49_U0.ap_done);
    assign proc_dep_vld_vec_25[3] = dl_detect_out ? proc_dep_vld_vec_25_reg[3] : (proc_25_data_FIFO_blk[3] | proc_25_data_PIPO_blk[3] | proc_25_start_FIFO_blk[3] | proc_25_TLF_FIFO_blk[3] | proc_25_input_sync_blk[3] | proc_25_output_sync_blk[3]);
    assign proc_25_data_FIFO_blk[4] = 1'b0;
    assign proc_25_data_PIPO_blk[4] = 1'b0;
    assign proc_25_start_FIFO_blk[4] = 1'b0;
    assign proc_25_TLF_FIFO_blk[4] = 1'b0;
    assign proc_25_input_sync_blk[4] = 1'b0;
    assign proc_25_output_sync_blk[4] = 1'b0 | (ap_done_reg_6 & write_back54_U0.ap_done & ~write_back50_U0.ap_done);
    assign proc_dep_vld_vec_25[4] = dl_detect_out ? proc_dep_vld_vec_25_reg[4] : (proc_25_data_FIFO_blk[4] | proc_25_data_PIPO_blk[4] | proc_25_start_FIFO_blk[4] | proc_25_TLF_FIFO_blk[4] | proc_25_input_sync_blk[4] | proc_25_output_sync_blk[4]);
    assign proc_25_data_FIFO_blk[5] = 1'b0;
    assign proc_25_data_PIPO_blk[5] = 1'b0;
    assign proc_25_start_FIFO_blk[5] = 1'b0;
    assign proc_25_TLF_FIFO_blk[5] = 1'b0;
    assign proc_25_input_sync_blk[5] = 1'b0;
    assign proc_25_output_sync_blk[5] = 1'b0 | (ap_done_reg_6 & write_back54_U0.ap_done & ~write_back51_U0.ap_done);
    assign proc_dep_vld_vec_25[5] = dl_detect_out ? proc_dep_vld_vec_25_reg[5] : (proc_25_data_FIFO_blk[5] | proc_25_data_PIPO_blk[5] | proc_25_start_FIFO_blk[5] | proc_25_TLF_FIFO_blk[5] | proc_25_input_sync_blk[5] | proc_25_output_sync_blk[5]);
    assign proc_25_data_FIFO_blk[6] = 1'b0;
    assign proc_25_data_PIPO_blk[6] = 1'b0;
    assign proc_25_start_FIFO_blk[6] = 1'b0;
    assign proc_25_TLF_FIFO_blk[6] = 1'b0;
    assign proc_25_input_sync_blk[6] = 1'b0;
    assign proc_25_output_sync_blk[6] = 1'b0 | (ap_done_reg_6 & write_back54_U0.ap_done & ~write_back52_U0.ap_done);
    assign proc_dep_vld_vec_25[6] = dl_detect_out ? proc_dep_vld_vec_25_reg[6] : (proc_25_data_FIFO_blk[6] | proc_25_data_PIPO_blk[6] | proc_25_start_FIFO_blk[6] | proc_25_TLF_FIFO_blk[6] | proc_25_input_sync_blk[6] | proc_25_output_sync_blk[6]);
    assign proc_25_data_FIFO_blk[7] = 1'b0;
    assign proc_25_data_PIPO_blk[7] = 1'b0;
    assign proc_25_start_FIFO_blk[7] = 1'b0;
    assign proc_25_TLF_FIFO_blk[7] = 1'b0;
    assign proc_25_input_sync_blk[7] = 1'b0;
    assign proc_25_output_sync_blk[7] = 1'b0 | (ap_done_reg_6 & write_back54_U0.ap_done & ~write_back53_U0.ap_done);
    assign proc_dep_vld_vec_25[7] = dl_detect_out ? proc_dep_vld_vec_25_reg[7] : (proc_25_data_FIFO_blk[7] | proc_25_data_PIPO_blk[7] | proc_25_start_FIFO_blk[7] | proc_25_TLF_FIFO_blk[7] | proc_25_input_sync_blk[7] | proc_25_output_sync_blk[7]);
    assign proc_25_data_FIFO_blk[8] = 1'b0;
    assign proc_25_data_PIPO_blk[8] = 1'b0;
    assign proc_25_start_FIFO_blk[8] = 1'b0;
    assign proc_25_TLF_FIFO_blk[8] = 1'b0;
    assign proc_25_input_sync_blk[8] = 1'b0;
    assign proc_25_output_sync_blk[8] = 1'b0 | (ap_done_reg_6 & write_back54_U0.ap_done & ~write_back55_U0.ap_done);
    assign proc_dep_vld_vec_25[8] = dl_detect_out ? proc_dep_vld_vec_25_reg[8] : (proc_25_data_FIFO_blk[8] | proc_25_data_PIPO_blk[8] | proc_25_start_FIFO_blk[8] | proc_25_TLF_FIFO_blk[8] | proc_25_input_sync_blk[8] | proc_25_output_sync_blk[8]);
    assign proc_25_data_FIFO_blk[9] = 1'b0;
    assign proc_25_data_PIPO_blk[9] = 1'b0;
    assign proc_25_start_FIFO_blk[9] = 1'b0;
    assign proc_25_TLF_FIFO_blk[9] = 1'b0;
    assign proc_25_input_sync_blk[9] = 1'b0;
    assign proc_25_output_sync_blk[9] = 1'b0 | (ap_done_reg_6 & write_back54_U0.ap_done & ~write_back56_U0.ap_done);
    assign proc_dep_vld_vec_25[9] = dl_detect_out ? proc_dep_vld_vec_25_reg[9] : (proc_25_data_FIFO_blk[9] | proc_25_data_PIPO_blk[9] | proc_25_start_FIFO_blk[9] | proc_25_TLF_FIFO_blk[9] | proc_25_input_sync_blk[9] | proc_25_output_sync_blk[9]);
    assign proc_25_data_FIFO_blk[10] = 1'b0;
    assign proc_25_data_PIPO_blk[10] = 1'b0;
    assign proc_25_start_FIFO_blk[10] = 1'b0;
    assign proc_25_TLF_FIFO_blk[10] = 1'b0;
    assign proc_25_input_sync_blk[10] = 1'b0;
    assign proc_25_output_sync_blk[10] = 1'b0 | (ap_done_reg_6 & write_back54_U0.ap_done & ~write_back57_U0.ap_done);
    assign proc_dep_vld_vec_25[10] = dl_detect_out ? proc_dep_vld_vec_25_reg[10] : (proc_25_data_FIFO_blk[10] | proc_25_data_PIPO_blk[10] | proc_25_start_FIFO_blk[10] | proc_25_TLF_FIFO_blk[10] | proc_25_input_sync_blk[10] | proc_25_output_sync_blk[10]);
    assign proc_25_data_FIFO_blk[11] = 1'b0;
    assign proc_25_data_PIPO_blk[11] = 1'b0;
    assign proc_25_start_FIFO_blk[11] = 1'b0;
    assign proc_25_TLF_FIFO_blk[11] = 1'b0;
    assign proc_25_input_sync_blk[11] = 1'b0;
    assign proc_25_output_sync_blk[11] = 1'b0 | (ap_done_reg_6 & write_back54_U0.ap_done & ~write_back58_U0.ap_done);
    assign proc_dep_vld_vec_25[11] = dl_detect_out ? proc_dep_vld_vec_25_reg[11] : (proc_25_data_FIFO_blk[11] | proc_25_data_PIPO_blk[11] | proc_25_start_FIFO_blk[11] | proc_25_TLF_FIFO_blk[11] | proc_25_input_sync_blk[11] | proc_25_output_sync_blk[11]);
    assign proc_25_data_FIFO_blk[12] = 1'b0;
    assign proc_25_data_PIPO_blk[12] = 1'b0;
    assign proc_25_start_FIFO_blk[12] = 1'b0;
    assign proc_25_TLF_FIFO_blk[12] = 1'b0;
    assign proc_25_input_sync_blk[12] = 1'b0;
    assign proc_25_output_sync_blk[12] = 1'b0 | (ap_done_reg_6 & write_back54_U0.ap_done & ~write_back59_U0.ap_done);
    assign proc_dep_vld_vec_25[12] = dl_detect_out ? proc_dep_vld_vec_25_reg[12] : (proc_25_data_FIFO_blk[12] | proc_25_data_PIPO_blk[12] | proc_25_start_FIFO_blk[12] | proc_25_TLF_FIFO_blk[12] | proc_25_input_sync_blk[12] | proc_25_output_sync_blk[12]);
    assign proc_25_data_FIFO_blk[13] = 1'b0;
    assign proc_25_data_PIPO_blk[13] = 1'b0;
    assign proc_25_start_FIFO_blk[13] = 1'b0;
    assign proc_25_TLF_FIFO_blk[13] = 1'b0;
    assign proc_25_input_sync_blk[13] = 1'b0;
    assign proc_25_output_sync_blk[13] = 1'b0 | (ap_done_reg_6 & write_back54_U0.ap_done & ~write_back60_U0.ap_done);
    assign proc_dep_vld_vec_25[13] = dl_detect_out ? proc_dep_vld_vec_25_reg[13] : (proc_25_data_FIFO_blk[13] | proc_25_data_PIPO_blk[13] | proc_25_start_FIFO_blk[13] | proc_25_TLF_FIFO_blk[13] | proc_25_input_sync_blk[13] | proc_25_output_sync_blk[13]);
    assign proc_25_data_FIFO_blk[14] = 1'b0;
    assign proc_25_data_PIPO_blk[14] = 1'b0;
    assign proc_25_start_FIFO_blk[14] = 1'b0;
    assign proc_25_TLF_FIFO_blk[14] = 1'b0;
    assign proc_25_input_sync_blk[14] = 1'b0;
    assign proc_25_output_sync_blk[14] = 1'b0 | (ap_done_reg_6 & write_back54_U0.ap_done & ~write_back61_U0.ap_done);
    assign proc_dep_vld_vec_25[14] = dl_detect_out ? proc_dep_vld_vec_25_reg[14] : (proc_25_data_FIFO_blk[14] | proc_25_data_PIPO_blk[14] | proc_25_start_FIFO_blk[14] | proc_25_TLF_FIFO_blk[14] | proc_25_input_sync_blk[14] | proc_25_output_sync_blk[14]);
    assign proc_25_data_FIFO_blk[15] = 1'b0;
    assign proc_25_data_PIPO_blk[15] = 1'b0;
    assign proc_25_start_FIFO_blk[15] = 1'b0;
    assign proc_25_TLF_FIFO_blk[15] = 1'b0;
    assign proc_25_input_sync_blk[15] = 1'b0;
    assign proc_25_output_sync_blk[15] = 1'b0 | (ap_done_reg_6 & write_back54_U0.ap_done & ~write_back62_U0.ap_done);
    assign proc_dep_vld_vec_25[15] = dl_detect_out ? proc_dep_vld_vec_25_reg[15] : (proc_25_data_FIFO_blk[15] | proc_25_data_PIPO_blk[15] | proc_25_start_FIFO_blk[15] | proc_25_TLF_FIFO_blk[15] | proc_25_input_sync_blk[15] | proc_25_output_sync_blk[15]);
    assign proc_25_data_FIFO_blk[16] = 1'b0;
    assign proc_25_data_PIPO_blk[16] = 1'b0;
    assign proc_25_start_FIFO_blk[16] = 1'b0;
    assign proc_25_TLF_FIFO_blk[16] = 1'b0;
    assign proc_25_input_sync_blk[16] = 1'b0;
    assign proc_25_output_sync_blk[16] = 1'b0 | (ap_done_reg_6 & write_back54_U0.ap_done & ~write_back63_U0.ap_done);
    assign proc_dep_vld_vec_25[16] = dl_detect_out ? proc_dep_vld_vec_25_reg[16] : (proc_25_data_FIFO_blk[16] | proc_25_data_PIPO_blk[16] | proc_25_start_FIFO_blk[16] | proc_25_TLF_FIFO_blk[16] | proc_25_input_sync_blk[16] | proc_25_output_sync_blk[16]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_25_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_25_reg <= proc_dep_vld_vec_25;
        end
    end
    assign in_chan_dep_vld_vec_25[0] = dep_chan_vld_0_25;
    assign in_chan_dep_data_vec_25[34 : 0] = dep_chan_data_0_25;
    assign token_in_vec_25[0] = token_0_25;
    assign in_chan_dep_vld_vec_25[1] = dep_chan_vld_9_25;
    assign in_chan_dep_data_vec_25[69 : 35] = dep_chan_data_9_25;
    assign token_in_vec_25[1] = token_9_25;
    assign in_chan_dep_vld_vec_25[2] = dep_chan_vld_19_25;
    assign in_chan_dep_data_vec_25[104 : 70] = dep_chan_data_19_25;
    assign token_in_vec_25[2] = token_19_25;
    assign in_chan_dep_vld_vec_25[3] = dep_chan_vld_20_25;
    assign in_chan_dep_data_vec_25[139 : 105] = dep_chan_data_20_25;
    assign token_in_vec_25[3] = token_20_25;
    assign in_chan_dep_vld_vec_25[4] = dep_chan_vld_21_25;
    assign in_chan_dep_data_vec_25[174 : 140] = dep_chan_data_21_25;
    assign token_in_vec_25[4] = token_21_25;
    assign in_chan_dep_vld_vec_25[5] = dep_chan_vld_22_25;
    assign in_chan_dep_data_vec_25[209 : 175] = dep_chan_data_22_25;
    assign token_in_vec_25[5] = token_22_25;
    assign in_chan_dep_vld_vec_25[6] = dep_chan_vld_23_25;
    assign in_chan_dep_data_vec_25[244 : 210] = dep_chan_data_23_25;
    assign token_in_vec_25[6] = token_23_25;
    assign in_chan_dep_vld_vec_25[7] = dep_chan_vld_24_25;
    assign in_chan_dep_data_vec_25[279 : 245] = dep_chan_data_24_25;
    assign token_in_vec_25[7] = token_24_25;
    assign in_chan_dep_vld_vec_25[8] = dep_chan_vld_26_25;
    assign in_chan_dep_data_vec_25[314 : 280] = dep_chan_data_26_25;
    assign token_in_vec_25[8] = token_26_25;
    assign in_chan_dep_vld_vec_25[9] = dep_chan_vld_27_25;
    assign in_chan_dep_data_vec_25[349 : 315] = dep_chan_data_27_25;
    assign token_in_vec_25[9] = token_27_25;
    assign in_chan_dep_vld_vec_25[10] = dep_chan_vld_28_25;
    assign in_chan_dep_data_vec_25[384 : 350] = dep_chan_data_28_25;
    assign token_in_vec_25[10] = token_28_25;
    assign in_chan_dep_vld_vec_25[11] = dep_chan_vld_29_25;
    assign in_chan_dep_data_vec_25[419 : 385] = dep_chan_data_29_25;
    assign token_in_vec_25[11] = token_29_25;
    assign in_chan_dep_vld_vec_25[12] = dep_chan_vld_30_25;
    assign in_chan_dep_data_vec_25[454 : 420] = dep_chan_data_30_25;
    assign token_in_vec_25[12] = token_30_25;
    assign in_chan_dep_vld_vec_25[13] = dep_chan_vld_31_25;
    assign in_chan_dep_data_vec_25[489 : 455] = dep_chan_data_31_25;
    assign token_in_vec_25[13] = token_31_25;
    assign in_chan_dep_vld_vec_25[14] = dep_chan_vld_32_25;
    assign in_chan_dep_data_vec_25[524 : 490] = dep_chan_data_32_25;
    assign token_in_vec_25[14] = token_32_25;
    assign in_chan_dep_vld_vec_25[15] = dep_chan_vld_33_25;
    assign in_chan_dep_data_vec_25[559 : 525] = dep_chan_data_33_25;
    assign token_in_vec_25[15] = token_33_25;
    assign in_chan_dep_vld_vec_25[16] = dep_chan_vld_34_25;
    assign in_chan_dep_data_vec_25[594 : 560] = dep_chan_data_34_25;
    assign token_in_vec_25[16] = token_34_25;
    assign dep_chan_vld_25_0 = out_chan_dep_vld_vec_25[0];
    assign dep_chan_data_25_0 = out_chan_dep_data_25;
    assign token_25_0 = token_out_vec_25[0];
    assign dep_chan_vld_25_9 = out_chan_dep_vld_vec_25[1];
    assign dep_chan_data_25_9 = out_chan_dep_data_25;
    assign token_25_9 = token_out_vec_25[1];
    assign dep_chan_vld_25_19 = out_chan_dep_vld_vec_25[2];
    assign dep_chan_data_25_19 = out_chan_dep_data_25;
    assign token_25_19 = token_out_vec_25[2];
    assign dep_chan_vld_25_20 = out_chan_dep_vld_vec_25[3];
    assign dep_chan_data_25_20 = out_chan_dep_data_25;
    assign token_25_20 = token_out_vec_25[3];
    assign dep_chan_vld_25_21 = out_chan_dep_vld_vec_25[4];
    assign dep_chan_data_25_21 = out_chan_dep_data_25;
    assign token_25_21 = token_out_vec_25[4];
    assign dep_chan_vld_25_22 = out_chan_dep_vld_vec_25[5];
    assign dep_chan_data_25_22 = out_chan_dep_data_25;
    assign token_25_22 = token_out_vec_25[5];
    assign dep_chan_vld_25_23 = out_chan_dep_vld_vec_25[6];
    assign dep_chan_data_25_23 = out_chan_dep_data_25;
    assign token_25_23 = token_out_vec_25[6];
    assign dep_chan_vld_25_24 = out_chan_dep_vld_vec_25[7];
    assign dep_chan_data_25_24 = out_chan_dep_data_25;
    assign token_25_24 = token_out_vec_25[7];
    assign dep_chan_vld_25_26 = out_chan_dep_vld_vec_25[8];
    assign dep_chan_data_25_26 = out_chan_dep_data_25;
    assign token_25_26 = token_out_vec_25[8];
    assign dep_chan_vld_25_27 = out_chan_dep_vld_vec_25[9];
    assign dep_chan_data_25_27 = out_chan_dep_data_25;
    assign token_25_27 = token_out_vec_25[9];
    assign dep_chan_vld_25_28 = out_chan_dep_vld_vec_25[10];
    assign dep_chan_data_25_28 = out_chan_dep_data_25;
    assign token_25_28 = token_out_vec_25[10];
    assign dep_chan_vld_25_29 = out_chan_dep_vld_vec_25[11];
    assign dep_chan_data_25_29 = out_chan_dep_data_25;
    assign token_25_29 = token_out_vec_25[11];
    assign dep_chan_vld_25_30 = out_chan_dep_vld_vec_25[12];
    assign dep_chan_data_25_30 = out_chan_dep_data_25;
    assign token_25_30 = token_out_vec_25[12];
    assign dep_chan_vld_25_31 = out_chan_dep_vld_vec_25[13];
    assign dep_chan_data_25_31 = out_chan_dep_data_25;
    assign token_25_31 = token_out_vec_25[13];
    assign dep_chan_vld_25_32 = out_chan_dep_vld_vec_25[14];
    assign dep_chan_data_25_32 = out_chan_dep_data_25;
    assign token_25_32 = token_out_vec_25[14];
    assign dep_chan_vld_25_33 = out_chan_dep_vld_vec_25[15];
    assign dep_chan_data_25_33 = out_chan_dep_data_25;
    assign token_25_33 = token_out_vec_25[15];
    assign dep_chan_vld_25_34 = out_chan_dep_vld_vec_25[16];
    assign dep_chan_data_25_34 = out_chan_dep_data_25;
    assign token_25_34 = token_out_vec_25[16];

    // Process: write_back55_U0
    kernel_pr_hls_deadlock_detect_unit #(35, 26, 17, 17) kernel_pr_hls_deadlock_detect_unit_26 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_26),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_26),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_26),
        .token_in_vec(token_in_vec_26),
        .dl_detect_in(dl_detect_out),
        .origin(origin[26]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_26),
        .out_chan_dep_data(out_chan_dep_data_26),
        .token_out_vec(token_out_vec_26),
        .dl_detect_out(dl_in_vec[26]));

    assign proc_26_data_FIFO_blk[0] = 1'b0 | (~write_back55_U0.H_blk_n) | (~write_back55_U0.hyperedge_size_blk_n);
    assign proc_26_data_PIPO_blk[0] = 1'b0;
    assign proc_26_start_FIFO_blk[0] = 1'b0 | (~start_for_write_back55_U0_U.if_empty_n & write_back55_U0.ap_idle & ~start_for_write_back55_U0_U.if_write);
    assign proc_26_TLF_FIFO_blk[0] = 1'b0;
    assign proc_26_input_sync_blk[0] = 1'b0;
    assign proc_26_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_26[0] = dl_detect_out ? proc_dep_vld_vec_26_reg[0] : (proc_26_data_FIFO_blk[0] | proc_26_data_PIPO_blk[0] | proc_26_start_FIFO_blk[0] | proc_26_TLF_FIFO_blk[0] | proc_26_input_sync_blk[0] | proc_26_output_sync_blk[0]);
    assign proc_26_data_FIFO_blk[1] = 1'b0 | (~write_back55_U0.value_stream_V_V7_blk_n);
    assign proc_26_data_PIPO_blk[1] = 1'b0;
    assign proc_26_start_FIFO_blk[1] = 1'b0;
    assign proc_26_TLF_FIFO_blk[1] = 1'b0;
    assign proc_26_input_sync_blk[1] = 1'b0;
    assign proc_26_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_26[1] = dl_detect_out ? proc_dep_vld_vec_26_reg[1] : (proc_26_data_FIFO_blk[1] | proc_26_data_PIPO_blk[1] | proc_26_start_FIFO_blk[1] | proc_26_TLF_FIFO_blk[1] | proc_26_input_sync_blk[1] | proc_26_output_sync_blk[1]);
    assign proc_26_data_FIFO_blk[2] = 1'b0;
    assign proc_26_data_PIPO_blk[2] = 1'b0;
    assign proc_26_start_FIFO_blk[2] = 1'b0;
    assign proc_26_TLF_FIFO_blk[2] = 1'b0;
    assign proc_26_input_sync_blk[2] = 1'b0;
    assign proc_26_output_sync_blk[2] = 1'b0 | (ap_done_reg_7 & write_back55_U0.ap_done & ~write_back48_U0.ap_done);
    assign proc_dep_vld_vec_26[2] = dl_detect_out ? proc_dep_vld_vec_26_reg[2] : (proc_26_data_FIFO_blk[2] | proc_26_data_PIPO_blk[2] | proc_26_start_FIFO_blk[2] | proc_26_TLF_FIFO_blk[2] | proc_26_input_sync_blk[2] | proc_26_output_sync_blk[2]);
    assign proc_26_data_FIFO_blk[3] = 1'b0;
    assign proc_26_data_PIPO_blk[3] = 1'b0;
    assign proc_26_start_FIFO_blk[3] = 1'b0;
    assign proc_26_TLF_FIFO_blk[3] = 1'b0;
    assign proc_26_input_sync_blk[3] = 1'b0;
    assign proc_26_output_sync_blk[3] = 1'b0 | (ap_done_reg_7 & write_back55_U0.ap_done & ~write_back49_U0.ap_done);
    assign proc_dep_vld_vec_26[3] = dl_detect_out ? proc_dep_vld_vec_26_reg[3] : (proc_26_data_FIFO_blk[3] | proc_26_data_PIPO_blk[3] | proc_26_start_FIFO_blk[3] | proc_26_TLF_FIFO_blk[3] | proc_26_input_sync_blk[3] | proc_26_output_sync_blk[3]);
    assign proc_26_data_FIFO_blk[4] = 1'b0;
    assign proc_26_data_PIPO_blk[4] = 1'b0;
    assign proc_26_start_FIFO_blk[4] = 1'b0;
    assign proc_26_TLF_FIFO_blk[4] = 1'b0;
    assign proc_26_input_sync_blk[4] = 1'b0;
    assign proc_26_output_sync_blk[4] = 1'b0 | (ap_done_reg_7 & write_back55_U0.ap_done & ~write_back50_U0.ap_done);
    assign proc_dep_vld_vec_26[4] = dl_detect_out ? proc_dep_vld_vec_26_reg[4] : (proc_26_data_FIFO_blk[4] | proc_26_data_PIPO_blk[4] | proc_26_start_FIFO_blk[4] | proc_26_TLF_FIFO_blk[4] | proc_26_input_sync_blk[4] | proc_26_output_sync_blk[4]);
    assign proc_26_data_FIFO_blk[5] = 1'b0;
    assign proc_26_data_PIPO_blk[5] = 1'b0;
    assign proc_26_start_FIFO_blk[5] = 1'b0;
    assign proc_26_TLF_FIFO_blk[5] = 1'b0;
    assign proc_26_input_sync_blk[5] = 1'b0;
    assign proc_26_output_sync_blk[5] = 1'b0 | (ap_done_reg_7 & write_back55_U0.ap_done & ~write_back51_U0.ap_done);
    assign proc_dep_vld_vec_26[5] = dl_detect_out ? proc_dep_vld_vec_26_reg[5] : (proc_26_data_FIFO_blk[5] | proc_26_data_PIPO_blk[5] | proc_26_start_FIFO_blk[5] | proc_26_TLF_FIFO_blk[5] | proc_26_input_sync_blk[5] | proc_26_output_sync_blk[5]);
    assign proc_26_data_FIFO_blk[6] = 1'b0;
    assign proc_26_data_PIPO_blk[6] = 1'b0;
    assign proc_26_start_FIFO_blk[6] = 1'b0;
    assign proc_26_TLF_FIFO_blk[6] = 1'b0;
    assign proc_26_input_sync_blk[6] = 1'b0;
    assign proc_26_output_sync_blk[6] = 1'b0 | (ap_done_reg_7 & write_back55_U0.ap_done & ~write_back52_U0.ap_done);
    assign proc_dep_vld_vec_26[6] = dl_detect_out ? proc_dep_vld_vec_26_reg[6] : (proc_26_data_FIFO_blk[6] | proc_26_data_PIPO_blk[6] | proc_26_start_FIFO_blk[6] | proc_26_TLF_FIFO_blk[6] | proc_26_input_sync_blk[6] | proc_26_output_sync_blk[6]);
    assign proc_26_data_FIFO_blk[7] = 1'b0;
    assign proc_26_data_PIPO_blk[7] = 1'b0;
    assign proc_26_start_FIFO_blk[7] = 1'b0;
    assign proc_26_TLF_FIFO_blk[7] = 1'b0;
    assign proc_26_input_sync_blk[7] = 1'b0;
    assign proc_26_output_sync_blk[7] = 1'b0 | (ap_done_reg_7 & write_back55_U0.ap_done & ~write_back53_U0.ap_done);
    assign proc_dep_vld_vec_26[7] = dl_detect_out ? proc_dep_vld_vec_26_reg[7] : (proc_26_data_FIFO_blk[7] | proc_26_data_PIPO_blk[7] | proc_26_start_FIFO_blk[7] | proc_26_TLF_FIFO_blk[7] | proc_26_input_sync_blk[7] | proc_26_output_sync_blk[7]);
    assign proc_26_data_FIFO_blk[8] = 1'b0;
    assign proc_26_data_PIPO_blk[8] = 1'b0;
    assign proc_26_start_FIFO_blk[8] = 1'b0;
    assign proc_26_TLF_FIFO_blk[8] = 1'b0;
    assign proc_26_input_sync_blk[8] = 1'b0;
    assign proc_26_output_sync_blk[8] = 1'b0 | (ap_done_reg_7 & write_back55_U0.ap_done & ~write_back54_U0.ap_done);
    assign proc_dep_vld_vec_26[8] = dl_detect_out ? proc_dep_vld_vec_26_reg[8] : (proc_26_data_FIFO_blk[8] | proc_26_data_PIPO_blk[8] | proc_26_start_FIFO_blk[8] | proc_26_TLF_FIFO_blk[8] | proc_26_input_sync_blk[8] | proc_26_output_sync_blk[8]);
    assign proc_26_data_FIFO_blk[9] = 1'b0;
    assign proc_26_data_PIPO_blk[9] = 1'b0;
    assign proc_26_start_FIFO_blk[9] = 1'b0;
    assign proc_26_TLF_FIFO_blk[9] = 1'b0;
    assign proc_26_input_sync_blk[9] = 1'b0;
    assign proc_26_output_sync_blk[9] = 1'b0 | (ap_done_reg_7 & write_back55_U0.ap_done & ~write_back56_U0.ap_done);
    assign proc_dep_vld_vec_26[9] = dl_detect_out ? proc_dep_vld_vec_26_reg[9] : (proc_26_data_FIFO_blk[9] | proc_26_data_PIPO_blk[9] | proc_26_start_FIFO_blk[9] | proc_26_TLF_FIFO_blk[9] | proc_26_input_sync_blk[9] | proc_26_output_sync_blk[9]);
    assign proc_26_data_FIFO_blk[10] = 1'b0;
    assign proc_26_data_PIPO_blk[10] = 1'b0;
    assign proc_26_start_FIFO_blk[10] = 1'b0;
    assign proc_26_TLF_FIFO_blk[10] = 1'b0;
    assign proc_26_input_sync_blk[10] = 1'b0;
    assign proc_26_output_sync_blk[10] = 1'b0 | (ap_done_reg_7 & write_back55_U0.ap_done & ~write_back57_U0.ap_done);
    assign proc_dep_vld_vec_26[10] = dl_detect_out ? proc_dep_vld_vec_26_reg[10] : (proc_26_data_FIFO_blk[10] | proc_26_data_PIPO_blk[10] | proc_26_start_FIFO_blk[10] | proc_26_TLF_FIFO_blk[10] | proc_26_input_sync_blk[10] | proc_26_output_sync_blk[10]);
    assign proc_26_data_FIFO_blk[11] = 1'b0;
    assign proc_26_data_PIPO_blk[11] = 1'b0;
    assign proc_26_start_FIFO_blk[11] = 1'b0;
    assign proc_26_TLF_FIFO_blk[11] = 1'b0;
    assign proc_26_input_sync_blk[11] = 1'b0;
    assign proc_26_output_sync_blk[11] = 1'b0 | (ap_done_reg_7 & write_back55_U0.ap_done & ~write_back58_U0.ap_done);
    assign proc_dep_vld_vec_26[11] = dl_detect_out ? proc_dep_vld_vec_26_reg[11] : (proc_26_data_FIFO_blk[11] | proc_26_data_PIPO_blk[11] | proc_26_start_FIFO_blk[11] | proc_26_TLF_FIFO_blk[11] | proc_26_input_sync_blk[11] | proc_26_output_sync_blk[11]);
    assign proc_26_data_FIFO_blk[12] = 1'b0;
    assign proc_26_data_PIPO_blk[12] = 1'b0;
    assign proc_26_start_FIFO_blk[12] = 1'b0;
    assign proc_26_TLF_FIFO_blk[12] = 1'b0;
    assign proc_26_input_sync_blk[12] = 1'b0;
    assign proc_26_output_sync_blk[12] = 1'b0 | (ap_done_reg_7 & write_back55_U0.ap_done & ~write_back59_U0.ap_done);
    assign proc_dep_vld_vec_26[12] = dl_detect_out ? proc_dep_vld_vec_26_reg[12] : (proc_26_data_FIFO_blk[12] | proc_26_data_PIPO_blk[12] | proc_26_start_FIFO_blk[12] | proc_26_TLF_FIFO_blk[12] | proc_26_input_sync_blk[12] | proc_26_output_sync_blk[12]);
    assign proc_26_data_FIFO_blk[13] = 1'b0;
    assign proc_26_data_PIPO_blk[13] = 1'b0;
    assign proc_26_start_FIFO_blk[13] = 1'b0;
    assign proc_26_TLF_FIFO_blk[13] = 1'b0;
    assign proc_26_input_sync_blk[13] = 1'b0;
    assign proc_26_output_sync_blk[13] = 1'b0 | (ap_done_reg_7 & write_back55_U0.ap_done & ~write_back60_U0.ap_done);
    assign proc_dep_vld_vec_26[13] = dl_detect_out ? proc_dep_vld_vec_26_reg[13] : (proc_26_data_FIFO_blk[13] | proc_26_data_PIPO_blk[13] | proc_26_start_FIFO_blk[13] | proc_26_TLF_FIFO_blk[13] | proc_26_input_sync_blk[13] | proc_26_output_sync_blk[13]);
    assign proc_26_data_FIFO_blk[14] = 1'b0;
    assign proc_26_data_PIPO_blk[14] = 1'b0;
    assign proc_26_start_FIFO_blk[14] = 1'b0;
    assign proc_26_TLF_FIFO_blk[14] = 1'b0;
    assign proc_26_input_sync_blk[14] = 1'b0;
    assign proc_26_output_sync_blk[14] = 1'b0 | (ap_done_reg_7 & write_back55_U0.ap_done & ~write_back61_U0.ap_done);
    assign proc_dep_vld_vec_26[14] = dl_detect_out ? proc_dep_vld_vec_26_reg[14] : (proc_26_data_FIFO_blk[14] | proc_26_data_PIPO_blk[14] | proc_26_start_FIFO_blk[14] | proc_26_TLF_FIFO_blk[14] | proc_26_input_sync_blk[14] | proc_26_output_sync_blk[14]);
    assign proc_26_data_FIFO_blk[15] = 1'b0;
    assign proc_26_data_PIPO_blk[15] = 1'b0;
    assign proc_26_start_FIFO_blk[15] = 1'b0;
    assign proc_26_TLF_FIFO_blk[15] = 1'b0;
    assign proc_26_input_sync_blk[15] = 1'b0;
    assign proc_26_output_sync_blk[15] = 1'b0 | (ap_done_reg_7 & write_back55_U0.ap_done & ~write_back62_U0.ap_done);
    assign proc_dep_vld_vec_26[15] = dl_detect_out ? proc_dep_vld_vec_26_reg[15] : (proc_26_data_FIFO_blk[15] | proc_26_data_PIPO_blk[15] | proc_26_start_FIFO_blk[15] | proc_26_TLF_FIFO_blk[15] | proc_26_input_sync_blk[15] | proc_26_output_sync_blk[15]);
    assign proc_26_data_FIFO_blk[16] = 1'b0;
    assign proc_26_data_PIPO_blk[16] = 1'b0;
    assign proc_26_start_FIFO_blk[16] = 1'b0;
    assign proc_26_TLF_FIFO_blk[16] = 1'b0;
    assign proc_26_input_sync_blk[16] = 1'b0;
    assign proc_26_output_sync_blk[16] = 1'b0 | (ap_done_reg_7 & write_back55_U0.ap_done & ~write_back63_U0.ap_done);
    assign proc_dep_vld_vec_26[16] = dl_detect_out ? proc_dep_vld_vec_26_reg[16] : (proc_26_data_FIFO_blk[16] | proc_26_data_PIPO_blk[16] | proc_26_start_FIFO_blk[16] | proc_26_TLF_FIFO_blk[16] | proc_26_input_sync_blk[16] | proc_26_output_sync_blk[16]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_26_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_26_reg <= proc_dep_vld_vec_26;
        end
    end
    assign in_chan_dep_vld_vec_26[0] = dep_chan_vld_0_26;
    assign in_chan_dep_data_vec_26[34 : 0] = dep_chan_data_0_26;
    assign token_in_vec_26[0] = token_0_26;
    assign in_chan_dep_vld_vec_26[1] = dep_chan_vld_10_26;
    assign in_chan_dep_data_vec_26[69 : 35] = dep_chan_data_10_26;
    assign token_in_vec_26[1] = token_10_26;
    assign in_chan_dep_vld_vec_26[2] = dep_chan_vld_19_26;
    assign in_chan_dep_data_vec_26[104 : 70] = dep_chan_data_19_26;
    assign token_in_vec_26[2] = token_19_26;
    assign in_chan_dep_vld_vec_26[3] = dep_chan_vld_20_26;
    assign in_chan_dep_data_vec_26[139 : 105] = dep_chan_data_20_26;
    assign token_in_vec_26[3] = token_20_26;
    assign in_chan_dep_vld_vec_26[4] = dep_chan_vld_21_26;
    assign in_chan_dep_data_vec_26[174 : 140] = dep_chan_data_21_26;
    assign token_in_vec_26[4] = token_21_26;
    assign in_chan_dep_vld_vec_26[5] = dep_chan_vld_22_26;
    assign in_chan_dep_data_vec_26[209 : 175] = dep_chan_data_22_26;
    assign token_in_vec_26[5] = token_22_26;
    assign in_chan_dep_vld_vec_26[6] = dep_chan_vld_23_26;
    assign in_chan_dep_data_vec_26[244 : 210] = dep_chan_data_23_26;
    assign token_in_vec_26[6] = token_23_26;
    assign in_chan_dep_vld_vec_26[7] = dep_chan_vld_24_26;
    assign in_chan_dep_data_vec_26[279 : 245] = dep_chan_data_24_26;
    assign token_in_vec_26[7] = token_24_26;
    assign in_chan_dep_vld_vec_26[8] = dep_chan_vld_25_26;
    assign in_chan_dep_data_vec_26[314 : 280] = dep_chan_data_25_26;
    assign token_in_vec_26[8] = token_25_26;
    assign in_chan_dep_vld_vec_26[9] = dep_chan_vld_27_26;
    assign in_chan_dep_data_vec_26[349 : 315] = dep_chan_data_27_26;
    assign token_in_vec_26[9] = token_27_26;
    assign in_chan_dep_vld_vec_26[10] = dep_chan_vld_28_26;
    assign in_chan_dep_data_vec_26[384 : 350] = dep_chan_data_28_26;
    assign token_in_vec_26[10] = token_28_26;
    assign in_chan_dep_vld_vec_26[11] = dep_chan_vld_29_26;
    assign in_chan_dep_data_vec_26[419 : 385] = dep_chan_data_29_26;
    assign token_in_vec_26[11] = token_29_26;
    assign in_chan_dep_vld_vec_26[12] = dep_chan_vld_30_26;
    assign in_chan_dep_data_vec_26[454 : 420] = dep_chan_data_30_26;
    assign token_in_vec_26[12] = token_30_26;
    assign in_chan_dep_vld_vec_26[13] = dep_chan_vld_31_26;
    assign in_chan_dep_data_vec_26[489 : 455] = dep_chan_data_31_26;
    assign token_in_vec_26[13] = token_31_26;
    assign in_chan_dep_vld_vec_26[14] = dep_chan_vld_32_26;
    assign in_chan_dep_data_vec_26[524 : 490] = dep_chan_data_32_26;
    assign token_in_vec_26[14] = token_32_26;
    assign in_chan_dep_vld_vec_26[15] = dep_chan_vld_33_26;
    assign in_chan_dep_data_vec_26[559 : 525] = dep_chan_data_33_26;
    assign token_in_vec_26[15] = token_33_26;
    assign in_chan_dep_vld_vec_26[16] = dep_chan_vld_34_26;
    assign in_chan_dep_data_vec_26[594 : 560] = dep_chan_data_34_26;
    assign token_in_vec_26[16] = token_34_26;
    assign dep_chan_vld_26_0 = out_chan_dep_vld_vec_26[0];
    assign dep_chan_data_26_0 = out_chan_dep_data_26;
    assign token_26_0 = token_out_vec_26[0];
    assign dep_chan_vld_26_10 = out_chan_dep_vld_vec_26[1];
    assign dep_chan_data_26_10 = out_chan_dep_data_26;
    assign token_26_10 = token_out_vec_26[1];
    assign dep_chan_vld_26_19 = out_chan_dep_vld_vec_26[2];
    assign dep_chan_data_26_19 = out_chan_dep_data_26;
    assign token_26_19 = token_out_vec_26[2];
    assign dep_chan_vld_26_20 = out_chan_dep_vld_vec_26[3];
    assign dep_chan_data_26_20 = out_chan_dep_data_26;
    assign token_26_20 = token_out_vec_26[3];
    assign dep_chan_vld_26_21 = out_chan_dep_vld_vec_26[4];
    assign dep_chan_data_26_21 = out_chan_dep_data_26;
    assign token_26_21 = token_out_vec_26[4];
    assign dep_chan_vld_26_22 = out_chan_dep_vld_vec_26[5];
    assign dep_chan_data_26_22 = out_chan_dep_data_26;
    assign token_26_22 = token_out_vec_26[5];
    assign dep_chan_vld_26_23 = out_chan_dep_vld_vec_26[6];
    assign dep_chan_data_26_23 = out_chan_dep_data_26;
    assign token_26_23 = token_out_vec_26[6];
    assign dep_chan_vld_26_24 = out_chan_dep_vld_vec_26[7];
    assign dep_chan_data_26_24 = out_chan_dep_data_26;
    assign token_26_24 = token_out_vec_26[7];
    assign dep_chan_vld_26_25 = out_chan_dep_vld_vec_26[8];
    assign dep_chan_data_26_25 = out_chan_dep_data_26;
    assign token_26_25 = token_out_vec_26[8];
    assign dep_chan_vld_26_27 = out_chan_dep_vld_vec_26[9];
    assign dep_chan_data_26_27 = out_chan_dep_data_26;
    assign token_26_27 = token_out_vec_26[9];
    assign dep_chan_vld_26_28 = out_chan_dep_vld_vec_26[10];
    assign dep_chan_data_26_28 = out_chan_dep_data_26;
    assign token_26_28 = token_out_vec_26[10];
    assign dep_chan_vld_26_29 = out_chan_dep_vld_vec_26[11];
    assign dep_chan_data_26_29 = out_chan_dep_data_26;
    assign token_26_29 = token_out_vec_26[11];
    assign dep_chan_vld_26_30 = out_chan_dep_vld_vec_26[12];
    assign dep_chan_data_26_30 = out_chan_dep_data_26;
    assign token_26_30 = token_out_vec_26[12];
    assign dep_chan_vld_26_31 = out_chan_dep_vld_vec_26[13];
    assign dep_chan_data_26_31 = out_chan_dep_data_26;
    assign token_26_31 = token_out_vec_26[13];
    assign dep_chan_vld_26_32 = out_chan_dep_vld_vec_26[14];
    assign dep_chan_data_26_32 = out_chan_dep_data_26;
    assign token_26_32 = token_out_vec_26[14];
    assign dep_chan_vld_26_33 = out_chan_dep_vld_vec_26[15];
    assign dep_chan_data_26_33 = out_chan_dep_data_26;
    assign token_26_33 = token_out_vec_26[15];
    assign dep_chan_vld_26_34 = out_chan_dep_vld_vec_26[16];
    assign dep_chan_data_26_34 = out_chan_dep_data_26;
    assign token_26_34 = token_out_vec_26[16];

    // Process: write_back56_U0
    kernel_pr_hls_deadlock_detect_unit #(35, 27, 17, 17) kernel_pr_hls_deadlock_detect_unit_27 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_27),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_27),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_27),
        .token_in_vec(token_in_vec_27),
        .dl_detect_in(dl_detect_out),
        .origin(origin[27]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_27),
        .out_chan_dep_data(out_chan_dep_data_27),
        .token_out_vec(token_out_vec_27),
        .dl_detect_out(dl_in_vec[27]));

    assign proc_27_data_FIFO_blk[0] = 1'b0 | (~write_back56_U0.H_blk_n) | (~write_back56_U0.hyperedge_size_blk_n);
    assign proc_27_data_PIPO_blk[0] = 1'b0;
    assign proc_27_start_FIFO_blk[0] = 1'b0 | (~start_for_write_back56_U0_U.if_empty_n & write_back56_U0.ap_idle & ~start_for_write_back56_U0_U.if_write);
    assign proc_27_TLF_FIFO_blk[0] = 1'b0;
    assign proc_27_input_sync_blk[0] = 1'b0;
    assign proc_27_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_27[0] = dl_detect_out ? proc_dep_vld_vec_27_reg[0] : (proc_27_data_FIFO_blk[0] | proc_27_data_PIPO_blk[0] | proc_27_start_FIFO_blk[0] | proc_27_TLF_FIFO_blk[0] | proc_27_input_sync_blk[0] | proc_27_output_sync_blk[0]);
    assign proc_27_data_FIFO_blk[1] = 1'b0 | (~write_back56_U0.value_stream_V_V8_blk_n);
    assign proc_27_data_PIPO_blk[1] = 1'b0;
    assign proc_27_start_FIFO_blk[1] = 1'b0;
    assign proc_27_TLF_FIFO_blk[1] = 1'b0;
    assign proc_27_input_sync_blk[1] = 1'b0;
    assign proc_27_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_27[1] = dl_detect_out ? proc_dep_vld_vec_27_reg[1] : (proc_27_data_FIFO_blk[1] | proc_27_data_PIPO_blk[1] | proc_27_start_FIFO_blk[1] | proc_27_TLF_FIFO_blk[1] | proc_27_input_sync_blk[1] | proc_27_output_sync_blk[1]);
    assign proc_27_data_FIFO_blk[2] = 1'b0;
    assign proc_27_data_PIPO_blk[2] = 1'b0;
    assign proc_27_start_FIFO_blk[2] = 1'b0;
    assign proc_27_TLF_FIFO_blk[2] = 1'b0;
    assign proc_27_input_sync_blk[2] = 1'b0;
    assign proc_27_output_sync_blk[2] = 1'b0 | (ap_done_reg_8 & write_back56_U0.ap_done & ~write_back48_U0.ap_done);
    assign proc_dep_vld_vec_27[2] = dl_detect_out ? proc_dep_vld_vec_27_reg[2] : (proc_27_data_FIFO_blk[2] | proc_27_data_PIPO_blk[2] | proc_27_start_FIFO_blk[2] | proc_27_TLF_FIFO_blk[2] | proc_27_input_sync_blk[2] | proc_27_output_sync_blk[2]);
    assign proc_27_data_FIFO_blk[3] = 1'b0;
    assign proc_27_data_PIPO_blk[3] = 1'b0;
    assign proc_27_start_FIFO_blk[3] = 1'b0;
    assign proc_27_TLF_FIFO_blk[3] = 1'b0;
    assign proc_27_input_sync_blk[3] = 1'b0;
    assign proc_27_output_sync_blk[3] = 1'b0 | (ap_done_reg_8 & write_back56_U0.ap_done & ~write_back49_U0.ap_done);
    assign proc_dep_vld_vec_27[3] = dl_detect_out ? proc_dep_vld_vec_27_reg[3] : (proc_27_data_FIFO_blk[3] | proc_27_data_PIPO_blk[3] | proc_27_start_FIFO_blk[3] | proc_27_TLF_FIFO_blk[3] | proc_27_input_sync_blk[3] | proc_27_output_sync_blk[3]);
    assign proc_27_data_FIFO_blk[4] = 1'b0;
    assign proc_27_data_PIPO_blk[4] = 1'b0;
    assign proc_27_start_FIFO_blk[4] = 1'b0;
    assign proc_27_TLF_FIFO_blk[4] = 1'b0;
    assign proc_27_input_sync_blk[4] = 1'b0;
    assign proc_27_output_sync_blk[4] = 1'b0 | (ap_done_reg_8 & write_back56_U0.ap_done & ~write_back50_U0.ap_done);
    assign proc_dep_vld_vec_27[4] = dl_detect_out ? proc_dep_vld_vec_27_reg[4] : (proc_27_data_FIFO_blk[4] | proc_27_data_PIPO_blk[4] | proc_27_start_FIFO_blk[4] | proc_27_TLF_FIFO_blk[4] | proc_27_input_sync_blk[4] | proc_27_output_sync_blk[4]);
    assign proc_27_data_FIFO_blk[5] = 1'b0;
    assign proc_27_data_PIPO_blk[5] = 1'b0;
    assign proc_27_start_FIFO_blk[5] = 1'b0;
    assign proc_27_TLF_FIFO_blk[5] = 1'b0;
    assign proc_27_input_sync_blk[5] = 1'b0;
    assign proc_27_output_sync_blk[5] = 1'b0 | (ap_done_reg_8 & write_back56_U0.ap_done & ~write_back51_U0.ap_done);
    assign proc_dep_vld_vec_27[5] = dl_detect_out ? proc_dep_vld_vec_27_reg[5] : (proc_27_data_FIFO_blk[5] | proc_27_data_PIPO_blk[5] | proc_27_start_FIFO_blk[5] | proc_27_TLF_FIFO_blk[5] | proc_27_input_sync_blk[5] | proc_27_output_sync_blk[5]);
    assign proc_27_data_FIFO_blk[6] = 1'b0;
    assign proc_27_data_PIPO_blk[6] = 1'b0;
    assign proc_27_start_FIFO_blk[6] = 1'b0;
    assign proc_27_TLF_FIFO_blk[6] = 1'b0;
    assign proc_27_input_sync_blk[6] = 1'b0;
    assign proc_27_output_sync_blk[6] = 1'b0 | (ap_done_reg_8 & write_back56_U0.ap_done & ~write_back52_U0.ap_done);
    assign proc_dep_vld_vec_27[6] = dl_detect_out ? proc_dep_vld_vec_27_reg[6] : (proc_27_data_FIFO_blk[6] | proc_27_data_PIPO_blk[6] | proc_27_start_FIFO_blk[6] | proc_27_TLF_FIFO_blk[6] | proc_27_input_sync_blk[6] | proc_27_output_sync_blk[6]);
    assign proc_27_data_FIFO_blk[7] = 1'b0;
    assign proc_27_data_PIPO_blk[7] = 1'b0;
    assign proc_27_start_FIFO_blk[7] = 1'b0;
    assign proc_27_TLF_FIFO_blk[7] = 1'b0;
    assign proc_27_input_sync_blk[7] = 1'b0;
    assign proc_27_output_sync_blk[7] = 1'b0 | (ap_done_reg_8 & write_back56_U0.ap_done & ~write_back53_U0.ap_done);
    assign proc_dep_vld_vec_27[7] = dl_detect_out ? proc_dep_vld_vec_27_reg[7] : (proc_27_data_FIFO_blk[7] | proc_27_data_PIPO_blk[7] | proc_27_start_FIFO_blk[7] | proc_27_TLF_FIFO_blk[7] | proc_27_input_sync_blk[7] | proc_27_output_sync_blk[7]);
    assign proc_27_data_FIFO_blk[8] = 1'b0;
    assign proc_27_data_PIPO_blk[8] = 1'b0;
    assign proc_27_start_FIFO_blk[8] = 1'b0;
    assign proc_27_TLF_FIFO_blk[8] = 1'b0;
    assign proc_27_input_sync_blk[8] = 1'b0;
    assign proc_27_output_sync_blk[8] = 1'b0 | (ap_done_reg_8 & write_back56_U0.ap_done & ~write_back54_U0.ap_done);
    assign proc_dep_vld_vec_27[8] = dl_detect_out ? proc_dep_vld_vec_27_reg[8] : (proc_27_data_FIFO_blk[8] | proc_27_data_PIPO_blk[8] | proc_27_start_FIFO_blk[8] | proc_27_TLF_FIFO_blk[8] | proc_27_input_sync_blk[8] | proc_27_output_sync_blk[8]);
    assign proc_27_data_FIFO_blk[9] = 1'b0;
    assign proc_27_data_PIPO_blk[9] = 1'b0;
    assign proc_27_start_FIFO_blk[9] = 1'b0;
    assign proc_27_TLF_FIFO_blk[9] = 1'b0;
    assign proc_27_input_sync_blk[9] = 1'b0;
    assign proc_27_output_sync_blk[9] = 1'b0 | (ap_done_reg_8 & write_back56_U0.ap_done & ~write_back55_U0.ap_done);
    assign proc_dep_vld_vec_27[9] = dl_detect_out ? proc_dep_vld_vec_27_reg[9] : (proc_27_data_FIFO_blk[9] | proc_27_data_PIPO_blk[9] | proc_27_start_FIFO_blk[9] | proc_27_TLF_FIFO_blk[9] | proc_27_input_sync_blk[9] | proc_27_output_sync_blk[9]);
    assign proc_27_data_FIFO_blk[10] = 1'b0;
    assign proc_27_data_PIPO_blk[10] = 1'b0;
    assign proc_27_start_FIFO_blk[10] = 1'b0;
    assign proc_27_TLF_FIFO_blk[10] = 1'b0;
    assign proc_27_input_sync_blk[10] = 1'b0;
    assign proc_27_output_sync_blk[10] = 1'b0 | (ap_done_reg_8 & write_back56_U0.ap_done & ~write_back57_U0.ap_done);
    assign proc_dep_vld_vec_27[10] = dl_detect_out ? proc_dep_vld_vec_27_reg[10] : (proc_27_data_FIFO_blk[10] | proc_27_data_PIPO_blk[10] | proc_27_start_FIFO_blk[10] | proc_27_TLF_FIFO_blk[10] | proc_27_input_sync_blk[10] | proc_27_output_sync_blk[10]);
    assign proc_27_data_FIFO_blk[11] = 1'b0;
    assign proc_27_data_PIPO_blk[11] = 1'b0;
    assign proc_27_start_FIFO_blk[11] = 1'b0;
    assign proc_27_TLF_FIFO_blk[11] = 1'b0;
    assign proc_27_input_sync_blk[11] = 1'b0;
    assign proc_27_output_sync_blk[11] = 1'b0 | (ap_done_reg_8 & write_back56_U0.ap_done & ~write_back58_U0.ap_done);
    assign proc_dep_vld_vec_27[11] = dl_detect_out ? proc_dep_vld_vec_27_reg[11] : (proc_27_data_FIFO_blk[11] | proc_27_data_PIPO_blk[11] | proc_27_start_FIFO_blk[11] | proc_27_TLF_FIFO_blk[11] | proc_27_input_sync_blk[11] | proc_27_output_sync_blk[11]);
    assign proc_27_data_FIFO_blk[12] = 1'b0;
    assign proc_27_data_PIPO_blk[12] = 1'b0;
    assign proc_27_start_FIFO_blk[12] = 1'b0;
    assign proc_27_TLF_FIFO_blk[12] = 1'b0;
    assign proc_27_input_sync_blk[12] = 1'b0;
    assign proc_27_output_sync_blk[12] = 1'b0 | (ap_done_reg_8 & write_back56_U0.ap_done & ~write_back59_U0.ap_done);
    assign proc_dep_vld_vec_27[12] = dl_detect_out ? proc_dep_vld_vec_27_reg[12] : (proc_27_data_FIFO_blk[12] | proc_27_data_PIPO_blk[12] | proc_27_start_FIFO_blk[12] | proc_27_TLF_FIFO_blk[12] | proc_27_input_sync_blk[12] | proc_27_output_sync_blk[12]);
    assign proc_27_data_FIFO_blk[13] = 1'b0;
    assign proc_27_data_PIPO_blk[13] = 1'b0;
    assign proc_27_start_FIFO_blk[13] = 1'b0;
    assign proc_27_TLF_FIFO_blk[13] = 1'b0;
    assign proc_27_input_sync_blk[13] = 1'b0;
    assign proc_27_output_sync_blk[13] = 1'b0 | (ap_done_reg_8 & write_back56_U0.ap_done & ~write_back60_U0.ap_done);
    assign proc_dep_vld_vec_27[13] = dl_detect_out ? proc_dep_vld_vec_27_reg[13] : (proc_27_data_FIFO_blk[13] | proc_27_data_PIPO_blk[13] | proc_27_start_FIFO_blk[13] | proc_27_TLF_FIFO_blk[13] | proc_27_input_sync_blk[13] | proc_27_output_sync_blk[13]);
    assign proc_27_data_FIFO_blk[14] = 1'b0;
    assign proc_27_data_PIPO_blk[14] = 1'b0;
    assign proc_27_start_FIFO_blk[14] = 1'b0;
    assign proc_27_TLF_FIFO_blk[14] = 1'b0;
    assign proc_27_input_sync_blk[14] = 1'b0;
    assign proc_27_output_sync_blk[14] = 1'b0 | (ap_done_reg_8 & write_back56_U0.ap_done & ~write_back61_U0.ap_done);
    assign proc_dep_vld_vec_27[14] = dl_detect_out ? proc_dep_vld_vec_27_reg[14] : (proc_27_data_FIFO_blk[14] | proc_27_data_PIPO_blk[14] | proc_27_start_FIFO_blk[14] | proc_27_TLF_FIFO_blk[14] | proc_27_input_sync_blk[14] | proc_27_output_sync_blk[14]);
    assign proc_27_data_FIFO_blk[15] = 1'b0;
    assign proc_27_data_PIPO_blk[15] = 1'b0;
    assign proc_27_start_FIFO_blk[15] = 1'b0;
    assign proc_27_TLF_FIFO_blk[15] = 1'b0;
    assign proc_27_input_sync_blk[15] = 1'b0;
    assign proc_27_output_sync_blk[15] = 1'b0 | (ap_done_reg_8 & write_back56_U0.ap_done & ~write_back62_U0.ap_done);
    assign proc_dep_vld_vec_27[15] = dl_detect_out ? proc_dep_vld_vec_27_reg[15] : (proc_27_data_FIFO_blk[15] | proc_27_data_PIPO_blk[15] | proc_27_start_FIFO_blk[15] | proc_27_TLF_FIFO_blk[15] | proc_27_input_sync_blk[15] | proc_27_output_sync_blk[15]);
    assign proc_27_data_FIFO_blk[16] = 1'b0;
    assign proc_27_data_PIPO_blk[16] = 1'b0;
    assign proc_27_start_FIFO_blk[16] = 1'b0;
    assign proc_27_TLF_FIFO_blk[16] = 1'b0;
    assign proc_27_input_sync_blk[16] = 1'b0;
    assign proc_27_output_sync_blk[16] = 1'b0 | (ap_done_reg_8 & write_back56_U0.ap_done & ~write_back63_U0.ap_done);
    assign proc_dep_vld_vec_27[16] = dl_detect_out ? proc_dep_vld_vec_27_reg[16] : (proc_27_data_FIFO_blk[16] | proc_27_data_PIPO_blk[16] | proc_27_start_FIFO_blk[16] | proc_27_TLF_FIFO_blk[16] | proc_27_input_sync_blk[16] | proc_27_output_sync_blk[16]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_27_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_27_reg <= proc_dep_vld_vec_27;
        end
    end
    assign in_chan_dep_vld_vec_27[0] = dep_chan_vld_0_27;
    assign in_chan_dep_data_vec_27[34 : 0] = dep_chan_data_0_27;
    assign token_in_vec_27[0] = token_0_27;
    assign in_chan_dep_vld_vec_27[1] = dep_chan_vld_11_27;
    assign in_chan_dep_data_vec_27[69 : 35] = dep_chan_data_11_27;
    assign token_in_vec_27[1] = token_11_27;
    assign in_chan_dep_vld_vec_27[2] = dep_chan_vld_19_27;
    assign in_chan_dep_data_vec_27[104 : 70] = dep_chan_data_19_27;
    assign token_in_vec_27[2] = token_19_27;
    assign in_chan_dep_vld_vec_27[3] = dep_chan_vld_20_27;
    assign in_chan_dep_data_vec_27[139 : 105] = dep_chan_data_20_27;
    assign token_in_vec_27[3] = token_20_27;
    assign in_chan_dep_vld_vec_27[4] = dep_chan_vld_21_27;
    assign in_chan_dep_data_vec_27[174 : 140] = dep_chan_data_21_27;
    assign token_in_vec_27[4] = token_21_27;
    assign in_chan_dep_vld_vec_27[5] = dep_chan_vld_22_27;
    assign in_chan_dep_data_vec_27[209 : 175] = dep_chan_data_22_27;
    assign token_in_vec_27[5] = token_22_27;
    assign in_chan_dep_vld_vec_27[6] = dep_chan_vld_23_27;
    assign in_chan_dep_data_vec_27[244 : 210] = dep_chan_data_23_27;
    assign token_in_vec_27[6] = token_23_27;
    assign in_chan_dep_vld_vec_27[7] = dep_chan_vld_24_27;
    assign in_chan_dep_data_vec_27[279 : 245] = dep_chan_data_24_27;
    assign token_in_vec_27[7] = token_24_27;
    assign in_chan_dep_vld_vec_27[8] = dep_chan_vld_25_27;
    assign in_chan_dep_data_vec_27[314 : 280] = dep_chan_data_25_27;
    assign token_in_vec_27[8] = token_25_27;
    assign in_chan_dep_vld_vec_27[9] = dep_chan_vld_26_27;
    assign in_chan_dep_data_vec_27[349 : 315] = dep_chan_data_26_27;
    assign token_in_vec_27[9] = token_26_27;
    assign in_chan_dep_vld_vec_27[10] = dep_chan_vld_28_27;
    assign in_chan_dep_data_vec_27[384 : 350] = dep_chan_data_28_27;
    assign token_in_vec_27[10] = token_28_27;
    assign in_chan_dep_vld_vec_27[11] = dep_chan_vld_29_27;
    assign in_chan_dep_data_vec_27[419 : 385] = dep_chan_data_29_27;
    assign token_in_vec_27[11] = token_29_27;
    assign in_chan_dep_vld_vec_27[12] = dep_chan_vld_30_27;
    assign in_chan_dep_data_vec_27[454 : 420] = dep_chan_data_30_27;
    assign token_in_vec_27[12] = token_30_27;
    assign in_chan_dep_vld_vec_27[13] = dep_chan_vld_31_27;
    assign in_chan_dep_data_vec_27[489 : 455] = dep_chan_data_31_27;
    assign token_in_vec_27[13] = token_31_27;
    assign in_chan_dep_vld_vec_27[14] = dep_chan_vld_32_27;
    assign in_chan_dep_data_vec_27[524 : 490] = dep_chan_data_32_27;
    assign token_in_vec_27[14] = token_32_27;
    assign in_chan_dep_vld_vec_27[15] = dep_chan_vld_33_27;
    assign in_chan_dep_data_vec_27[559 : 525] = dep_chan_data_33_27;
    assign token_in_vec_27[15] = token_33_27;
    assign in_chan_dep_vld_vec_27[16] = dep_chan_vld_34_27;
    assign in_chan_dep_data_vec_27[594 : 560] = dep_chan_data_34_27;
    assign token_in_vec_27[16] = token_34_27;
    assign dep_chan_vld_27_0 = out_chan_dep_vld_vec_27[0];
    assign dep_chan_data_27_0 = out_chan_dep_data_27;
    assign token_27_0 = token_out_vec_27[0];
    assign dep_chan_vld_27_11 = out_chan_dep_vld_vec_27[1];
    assign dep_chan_data_27_11 = out_chan_dep_data_27;
    assign token_27_11 = token_out_vec_27[1];
    assign dep_chan_vld_27_19 = out_chan_dep_vld_vec_27[2];
    assign dep_chan_data_27_19 = out_chan_dep_data_27;
    assign token_27_19 = token_out_vec_27[2];
    assign dep_chan_vld_27_20 = out_chan_dep_vld_vec_27[3];
    assign dep_chan_data_27_20 = out_chan_dep_data_27;
    assign token_27_20 = token_out_vec_27[3];
    assign dep_chan_vld_27_21 = out_chan_dep_vld_vec_27[4];
    assign dep_chan_data_27_21 = out_chan_dep_data_27;
    assign token_27_21 = token_out_vec_27[4];
    assign dep_chan_vld_27_22 = out_chan_dep_vld_vec_27[5];
    assign dep_chan_data_27_22 = out_chan_dep_data_27;
    assign token_27_22 = token_out_vec_27[5];
    assign dep_chan_vld_27_23 = out_chan_dep_vld_vec_27[6];
    assign dep_chan_data_27_23 = out_chan_dep_data_27;
    assign token_27_23 = token_out_vec_27[6];
    assign dep_chan_vld_27_24 = out_chan_dep_vld_vec_27[7];
    assign dep_chan_data_27_24 = out_chan_dep_data_27;
    assign token_27_24 = token_out_vec_27[7];
    assign dep_chan_vld_27_25 = out_chan_dep_vld_vec_27[8];
    assign dep_chan_data_27_25 = out_chan_dep_data_27;
    assign token_27_25 = token_out_vec_27[8];
    assign dep_chan_vld_27_26 = out_chan_dep_vld_vec_27[9];
    assign dep_chan_data_27_26 = out_chan_dep_data_27;
    assign token_27_26 = token_out_vec_27[9];
    assign dep_chan_vld_27_28 = out_chan_dep_vld_vec_27[10];
    assign dep_chan_data_27_28 = out_chan_dep_data_27;
    assign token_27_28 = token_out_vec_27[10];
    assign dep_chan_vld_27_29 = out_chan_dep_vld_vec_27[11];
    assign dep_chan_data_27_29 = out_chan_dep_data_27;
    assign token_27_29 = token_out_vec_27[11];
    assign dep_chan_vld_27_30 = out_chan_dep_vld_vec_27[12];
    assign dep_chan_data_27_30 = out_chan_dep_data_27;
    assign token_27_30 = token_out_vec_27[12];
    assign dep_chan_vld_27_31 = out_chan_dep_vld_vec_27[13];
    assign dep_chan_data_27_31 = out_chan_dep_data_27;
    assign token_27_31 = token_out_vec_27[13];
    assign dep_chan_vld_27_32 = out_chan_dep_vld_vec_27[14];
    assign dep_chan_data_27_32 = out_chan_dep_data_27;
    assign token_27_32 = token_out_vec_27[14];
    assign dep_chan_vld_27_33 = out_chan_dep_vld_vec_27[15];
    assign dep_chan_data_27_33 = out_chan_dep_data_27;
    assign token_27_33 = token_out_vec_27[15];
    assign dep_chan_vld_27_34 = out_chan_dep_vld_vec_27[16];
    assign dep_chan_data_27_34 = out_chan_dep_data_27;
    assign token_27_34 = token_out_vec_27[16];

    // Process: write_back57_U0
    kernel_pr_hls_deadlock_detect_unit #(35, 28, 17, 17) kernel_pr_hls_deadlock_detect_unit_28 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_28),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_28),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_28),
        .token_in_vec(token_in_vec_28),
        .dl_detect_in(dl_detect_out),
        .origin(origin[28]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_28),
        .out_chan_dep_data(out_chan_dep_data_28),
        .token_out_vec(token_out_vec_28),
        .dl_detect_out(dl_in_vec[28]));

    assign proc_28_data_FIFO_blk[0] = 1'b0 | (~write_back57_U0.H_blk_n) | (~write_back57_U0.hyperedge_size_blk_n);
    assign proc_28_data_PIPO_blk[0] = 1'b0;
    assign proc_28_start_FIFO_blk[0] = 1'b0 | (~start_for_write_back57_U0_U.if_empty_n & write_back57_U0.ap_idle & ~start_for_write_back57_U0_U.if_write);
    assign proc_28_TLF_FIFO_blk[0] = 1'b0;
    assign proc_28_input_sync_blk[0] = 1'b0;
    assign proc_28_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_28[0] = dl_detect_out ? proc_dep_vld_vec_28_reg[0] : (proc_28_data_FIFO_blk[0] | proc_28_data_PIPO_blk[0] | proc_28_start_FIFO_blk[0] | proc_28_TLF_FIFO_blk[0] | proc_28_input_sync_blk[0] | proc_28_output_sync_blk[0]);
    assign proc_28_data_FIFO_blk[1] = 1'b0 | (~write_back57_U0.value_stream_V_V9_blk_n);
    assign proc_28_data_PIPO_blk[1] = 1'b0;
    assign proc_28_start_FIFO_blk[1] = 1'b0;
    assign proc_28_TLF_FIFO_blk[1] = 1'b0;
    assign proc_28_input_sync_blk[1] = 1'b0;
    assign proc_28_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_28[1] = dl_detect_out ? proc_dep_vld_vec_28_reg[1] : (proc_28_data_FIFO_blk[1] | proc_28_data_PIPO_blk[1] | proc_28_start_FIFO_blk[1] | proc_28_TLF_FIFO_blk[1] | proc_28_input_sync_blk[1] | proc_28_output_sync_blk[1]);
    assign proc_28_data_FIFO_blk[2] = 1'b0;
    assign proc_28_data_PIPO_blk[2] = 1'b0;
    assign proc_28_start_FIFO_blk[2] = 1'b0;
    assign proc_28_TLF_FIFO_blk[2] = 1'b0;
    assign proc_28_input_sync_blk[2] = 1'b0;
    assign proc_28_output_sync_blk[2] = 1'b0 | (ap_done_reg_9 & write_back57_U0.ap_done & ~write_back48_U0.ap_done);
    assign proc_dep_vld_vec_28[2] = dl_detect_out ? proc_dep_vld_vec_28_reg[2] : (proc_28_data_FIFO_blk[2] | proc_28_data_PIPO_blk[2] | proc_28_start_FIFO_blk[2] | proc_28_TLF_FIFO_blk[2] | proc_28_input_sync_blk[2] | proc_28_output_sync_blk[2]);
    assign proc_28_data_FIFO_blk[3] = 1'b0;
    assign proc_28_data_PIPO_blk[3] = 1'b0;
    assign proc_28_start_FIFO_blk[3] = 1'b0;
    assign proc_28_TLF_FIFO_blk[3] = 1'b0;
    assign proc_28_input_sync_blk[3] = 1'b0;
    assign proc_28_output_sync_blk[3] = 1'b0 | (ap_done_reg_9 & write_back57_U0.ap_done & ~write_back49_U0.ap_done);
    assign proc_dep_vld_vec_28[3] = dl_detect_out ? proc_dep_vld_vec_28_reg[3] : (proc_28_data_FIFO_blk[3] | proc_28_data_PIPO_blk[3] | proc_28_start_FIFO_blk[3] | proc_28_TLF_FIFO_blk[3] | proc_28_input_sync_blk[3] | proc_28_output_sync_blk[3]);
    assign proc_28_data_FIFO_blk[4] = 1'b0;
    assign proc_28_data_PIPO_blk[4] = 1'b0;
    assign proc_28_start_FIFO_blk[4] = 1'b0;
    assign proc_28_TLF_FIFO_blk[4] = 1'b0;
    assign proc_28_input_sync_blk[4] = 1'b0;
    assign proc_28_output_sync_blk[4] = 1'b0 | (ap_done_reg_9 & write_back57_U0.ap_done & ~write_back50_U0.ap_done);
    assign proc_dep_vld_vec_28[4] = dl_detect_out ? proc_dep_vld_vec_28_reg[4] : (proc_28_data_FIFO_blk[4] | proc_28_data_PIPO_blk[4] | proc_28_start_FIFO_blk[4] | proc_28_TLF_FIFO_blk[4] | proc_28_input_sync_blk[4] | proc_28_output_sync_blk[4]);
    assign proc_28_data_FIFO_blk[5] = 1'b0;
    assign proc_28_data_PIPO_blk[5] = 1'b0;
    assign proc_28_start_FIFO_blk[5] = 1'b0;
    assign proc_28_TLF_FIFO_blk[5] = 1'b0;
    assign proc_28_input_sync_blk[5] = 1'b0;
    assign proc_28_output_sync_blk[5] = 1'b0 | (ap_done_reg_9 & write_back57_U0.ap_done & ~write_back51_U0.ap_done);
    assign proc_dep_vld_vec_28[5] = dl_detect_out ? proc_dep_vld_vec_28_reg[5] : (proc_28_data_FIFO_blk[5] | proc_28_data_PIPO_blk[5] | proc_28_start_FIFO_blk[5] | proc_28_TLF_FIFO_blk[5] | proc_28_input_sync_blk[5] | proc_28_output_sync_blk[5]);
    assign proc_28_data_FIFO_blk[6] = 1'b0;
    assign proc_28_data_PIPO_blk[6] = 1'b0;
    assign proc_28_start_FIFO_blk[6] = 1'b0;
    assign proc_28_TLF_FIFO_blk[6] = 1'b0;
    assign proc_28_input_sync_blk[6] = 1'b0;
    assign proc_28_output_sync_blk[6] = 1'b0 | (ap_done_reg_9 & write_back57_U0.ap_done & ~write_back52_U0.ap_done);
    assign proc_dep_vld_vec_28[6] = dl_detect_out ? proc_dep_vld_vec_28_reg[6] : (proc_28_data_FIFO_blk[6] | proc_28_data_PIPO_blk[6] | proc_28_start_FIFO_blk[6] | proc_28_TLF_FIFO_blk[6] | proc_28_input_sync_blk[6] | proc_28_output_sync_blk[6]);
    assign proc_28_data_FIFO_blk[7] = 1'b0;
    assign proc_28_data_PIPO_blk[7] = 1'b0;
    assign proc_28_start_FIFO_blk[7] = 1'b0;
    assign proc_28_TLF_FIFO_blk[7] = 1'b0;
    assign proc_28_input_sync_blk[7] = 1'b0;
    assign proc_28_output_sync_blk[7] = 1'b0 | (ap_done_reg_9 & write_back57_U0.ap_done & ~write_back53_U0.ap_done);
    assign proc_dep_vld_vec_28[7] = dl_detect_out ? proc_dep_vld_vec_28_reg[7] : (proc_28_data_FIFO_blk[7] | proc_28_data_PIPO_blk[7] | proc_28_start_FIFO_blk[7] | proc_28_TLF_FIFO_blk[7] | proc_28_input_sync_blk[7] | proc_28_output_sync_blk[7]);
    assign proc_28_data_FIFO_blk[8] = 1'b0;
    assign proc_28_data_PIPO_blk[8] = 1'b0;
    assign proc_28_start_FIFO_blk[8] = 1'b0;
    assign proc_28_TLF_FIFO_blk[8] = 1'b0;
    assign proc_28_input_sync_blk[8] = 1'b0;
    assign proc_28_output_sync_blk[8] = 1'b0 | (ap_done_reg_9 & write_back57_U0.ap_done & ~write_back54_U0.ap_done);
    assign proc_dep_vld_vec_28[8] = dl_detect_out ? proc_dep_vld_vec_28_reg[8] : (proc_28_data_FIFO_blk[8] | proc_28_data_PIPO_blk[8] | proc_28_start_FIFO_blk[8] | proc_28_TLF_FIFO_blk[8] | proc_28_input_sync_blk[8] | proc_28_output_sync_blk[8]);
    assign proc_28_data_FIFO_blk[9] = 1'b0;
    assign proc_28_data_PIPO_blk[9] = 1'b0;
    assign proc_28_start_FIFO_blk[9] = 1'b0;
    assign proc_28_TLF_FIFO_blk[9] = 1'b0;
    assign proc_28_input_sync_blk[9] = 1'b0;
    assign proc_28_output_sync_blk[9] = 1'b0 | (ap_done_reg_9 & write_back57_U0.ap_done & ~write_back55_U0.ap_done);
    assign proc_dep_vld_vec_28[9] = dl_detect_out ? proc_dep_vld_vec_28_reg[9] : (proc_28_data_FIFO_blk[9] | proc_28_data_PIPO_blk[9] | proc_28_start_FIFO_blk[9] | proc_28_TLF_FIFO_blk[9] | proc_28_input_sync_blk[9] | proc_28_output_sync_blk[9]);
    assign proc_28_data_FIFO_blk[10] = 1'b0;
    assign proc_28_data_PIPO_blk[10] = 1'b0;
    assign proc_28_start_FIFO_blk[10] = 1'b0;
    assign proc_28_TLF_FIFO_blk[10] = 1'b0;
    assign proc_28_input_sync_blk[10] = 1'b0;
    assign proc_28_output_sync_blk[10] = 1'b0 | (ap_done_reg_9 & write_back57_U0.ap_done & ~write_back56_U0.ap_done);
    assign proc_dep_vld_vec_28[10] = dl_detect_out ? proc_dep_vld_vec_28_reg[10] : (proc_28_data_FIFO_blk[10] | proc_28_data_PIPO_blk[10] | proc_28_start_FIFO_blk[10] | proc_28_TLF_FIFO_blk[10] | proc_28_input_sync_blk[10] | proc_28_output_sync_blk[10]);
    assign proc_28_data_FIFO_blk[11] = 1'b0;
    assign proc_28_data_PIPO_blk[11] = 1'b0;
    assign proc_28_start_FIFO_blk[11] = 1'b0;
    assign proc_28_TLF_FIFO_blk[11] = 1'b0;
    assign proc_28_input_sync_blk[11] = 1'b0;
    assign proc_28_output_sync_blk[11] = 1'b0 | (ap_done_reg_9 & write_back57_U0.ap_done & ~write_back58_U0.ap_done);
    assign proc_dep_vld_vec_28[11] = dl_detect_out ? proc_dep_vld_vec_28_reg[11] : (proc_28_data_FIFO_blk[11] | proc_28_data_PIPO_blk[11] | proc_28_start_FIFO_blk[11] | proc_28_TLF_FIFO_blk[11] | proc_28_input_sync_blk[11] | proc_28_output_sync_blk[11]);
    assign proc_28_data_FIFO_blk[12] = 1'b0;
    assign proc_28_data_PIPO_blk[12] = 1'b0;
    assign proc_28_start_FIFO_blk[12] = 1'b0;
    assign proc_28_TLF_FIFO_blk[12] = 1'b0;
    assign proc_28_input_sync_blk[12] = 1'b0;
    assign proc_28_output_sync_blk[12] = 1'b0 | (ap_done_reg_9 & write_back57_U0.ap_done & ~write_back59_U0.ap_done);
    assign proc_dep_vld_vec_28[12] = dl_detect_out ? proc_dep_vld_vec_28_reg[12] : (proc_28_data_FIFO_blk[12] | proc_28_data_PIPO_blk[12] | proc_28_start_FIFO_blk[12] | proc_28_TLF_FIFO_blk[12] | proc_28_input_sync_blk[12] | proc_28_output_sync_blk[12]);
    assign proc_28_data_FIFO_blk[13] = 1'b0;
    assign proc_28_data_PIPO_blk[13] = 1'b0;
    assign proc_28_start_FIFO_blk[13] = 1'b0;
    assign proc_28_TLF_FIFO_blk[13] = 1'b0;
    assign proc_28_input_sync_blk[13] = 1'b0;
    assign proc_28_output_sync_blk[13] = 1'b0 | (ap_done_reg_9 & write_back57_U0.ap_done & ~write_back60_U0.ap_done);
    assign proc_dep_vld_vec_28[13] = dl_detect_out ? proc_dep_vld_vec_28_reg[13] : (proc_28_data_FIFO_blk[13] | proc_28_data_PIPO_blk[13] | proc_28_start_FIFO_blk[13] | proc_28_TLF_FIFO_blk[13] | proc_28_input_sync_blk[13] | proc_28_output_sync_blk[13]);
    assign proc_28_data_FIFO_blk[14] = 1'b0;
    assign proc_28_data_PIPO_blk[14] = 1'b0;
    assign proc_28_start_FIFO_blk[14] = 1'b0;
    assign proc_28_TLF_FIFO_blk[14] = 1'b0;
    assign proc_28_input_sync_blk[14] = 1'b0;
    assign proc_28_output_sync_blk[14] = 1'b0 | (ap_done_reg_9 & write_back57_U0.ap_done & ~write_back61_U0.ap_done);
    assign proc_dep_vld_vec_28[14] = dl_detect_out ? proc_dep_vld_vec_28_reg[14] : (proc_28_data_FIFO_blk[14] | proc_28_data_PIPO_blk[14] | proc_28_start_FIFO_blk[14] | proc_28_TLF_FIFO_blk[14] | proc_28_input_sync_blk[14] | proc_28_output_sync_blk[14]);
    assign proc_28_data_FIFO_blk[15] = 1'b0;
    assign proc_28_data_PIPO_blk[15] = 1'b0;
    assign proc_28_start_FIFO_blk[15] = 1'b0;
    assign proc_28_TLF_FIFO_blk[15] = 1'b0;
    assign proc_28_input_sync_blk[15] = 1'b0;
    assign proc_28_output_sync_blk[15] = 1'b0 | (ap_done_reg_9 & write_back57_U0.ap_done & ~write_back62_U0.ap_done);
    assign proc_dep_vld_vec_28[15] = dl_detect_out ? proc_dep_vld_vec_28_reg[15] : (proc_28_data_FIFO_blk[15] | proc_28_data_PIPO_blk[15] | proc_28_start_FIFO_blk[15] | proc_28_TLF_FIFO_blk[15] | proc_28_input_sync_blk[15] | proc_28_output_sync_blk[15]);
    assign proc_28_data_FIFO_blk[16] = 1'b0;
    assign proc_28_data_PIPO_blk[16] = 1'b0;
    assign proc_28_start_FIFO_blk[16] = 1'b0;
    assign proc_28_TLF_FIFO_blk[16] = 1'b0;
    assign proc_28_input_sync_blk[16] = 1'b0;
    assign proc_28_output_sync_blk[16] = 1'b0 | (ap_done_reg_9 & write_back57_U0.ap_done & ~write_back63_U0.ap_done);
    assign proc_dep_vld_vec_28[16] = dl_detect_out ? proc_dep_vld_vec_28_reg[16] : (proc_28_data_FIFO_blk[16] | proc_28_data_PIPO_blk[16] | proc_28_start_FIFO_blk[16] | proc_28_TLF_FIFO_blk[16] | proc_28_input_sync_blk[16] | proc_28_output_sync_blk[16]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_28_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_28_reg <= proc_dep_vld_vec_28;
        end
    end
    assign in_chan_dep_vld_vec_28[0] = dep_chan_vld_0_28;
    assign in_chan_dep_data_vec_28[34 : 0] = dep_chan_data_0_28;
    assign token_in_vec_28[0] = token_0_28;
    assign in_chan_dep_vld_vec_28[1] = dep_chan_vld_12_28;
    assign in_chan_dep_data_vec_28[69 : 35] = dep_chan_data_12_28;
    assign token_in_vec_28[1] = token_12_28;
    assign in_chan_dep_vld_vec_28[2] = dep_chan_vld_19_28;
    assign in_chan_dep_data_vec_28[104 : 70] = dep_chan_data_19_28;
    assign token_in_vec_28[2] = token_19_28;
    assign in_chan_dep_vld_vec_28[3] = dep_chan_vld_20_28;
    assign in_chan_dep_data_vec_28[139 : 105] = dep_chan_data_20_28;
    assign token_in_vec_28[3] = token_20_28;
    assign in_chan_dep_vld_vec_28[4] = dep_chan_vld_21_28;
    assign in_chan_dep_data_vec_28[174 : 140] = dep_chan_data_21_28;
    assign token_in_vec_28[4] = token_21_28;
    assign in_chan_dep_vld_vec_28[5] = dep_chan_vld_22_28;
    assign in_chan_dep_data_vec_28[209 : 175] = dep_chan_data_22_28;
    assign token_in_vec_28[5] = token_22_28;
    assign in_chan_dep_vld_vec_28[6] = dep_chan_vld_23_28;
    assign in_chan_dep_data_vec_28[244 : 210] = dep_chan_data_23_28;
    assign token_in_vec_28[6] = token_23_28;
    assign in_chan_dep_vld_vec_28[7] = dep_chan_vld_24_28;
    assign in_chan_dep_data_vec_28[279 : 245] = dep_chan_data_24_28;
    assign token_in_vec_28[7] = token_24_28;
    assign in_chan_dep_vld_vec_28[8] = dep_chan_vld_25_28;
    assign in_chan_dep_data_vec_28[314 : 280] = dep_chan_data_25_28;
    assign token_in_vec_28[8] = token_25_28;
    assign in_chan_dep_vld_vec_28[9] = dep_chan_vld_26_28;
    assign in_chan_dep_data_vec_28[349 : 315] = dep_chan_data_26_28;
    assign token_in_vec_28[9] = token_26_28;
    assign in_chan_dep_vld_vec_28[10] = dep_chan_vld_27_28;
    assign in_chan_dep_data_vec_28[384 : 350] = dep_chan_data_27_28;
    assign token_in_vec_28[10] = token_27_28;
    assign in_chan_dep_vld_vec_28[11] = dep_chan_vld_29_28;
    assign in_chan_dep_data_vec_28[419 : 385] = dep_chan_data_29_28;
    assign token_in_vec_28[11] = token_29_28;
    assign in_chan_dep_vld_vec_28[12] = dep_chan_vld_30_28;
    assign in_chan_dep_data_vec_28[454 : 420] = dep_chan_data_30_28;
    assign token_in_vec_28[12] = token_30_28;
    assign in_chan_dep_vld_vec_28[13] = dep_chan_vld_31_28;
    assign in_chan_dep_data_vec_28[489 : 455] = dep_chan_data_31_28;
    assign token_in_vec_28[13] = token_31_28;
    assign in_chan_dep_vld_vec_28[14] = dep_chan_vld_32_28;
    assign in_chan_dep_data_vec_28[524 : 490] = dep_chan_data_32_28;
    assign token_in_vec_28[14] = token_32_28;
    assign in_chan_dep_vld_vec_28[15] = dep_chan_vld_33_28;
    assign in_chan_dep_data_vec_28[559 : 525] = dep_chan_data_33_28;
    assign token_in_vec_28[15] = token_33_28;
    assign in_chan_dep_vld_vec_28[16] = dep_chan_vld_34_28;
    assign in_chan_dep_data_vec_28[594 : 560] = dep_chan_data_34_28;
    assign token_in_vec_28[16] = token_34_28;
    assign dep_chan_vld_28_0 = out_chan_dep_vld_vec_28[0];
    assign dep_chan_data_28_0 = out_chan_dep_data_28;
    assign token_28_0 = token_out_vec_28[0];
    assign dep_chan_vld_28_12 = out_chan_dep_vld_vec_28[1];
    assign dep_chan_data_28_12 = out_chan_dep_data_28;
    assign token_28_12 = token_out_vec_28[1];
    assign dep_chan_vld_28_19 = out_chan_dep_vld_vec_28[2];
    assign dep_chan_data_28_19 = out_chan_dep_data_28;
    assign token_28_19 = token_out_vec_28[2];
    assign dep_chan_vld_28_20 = out_chan_dep_vld_vec_28[3];
    assign dep_chan_data_28_20 = out_chan_dep_data_28;
    assign token_28_20 = token_out_vec_28[3];
    assign dep_chan_vld_28_21 = out_chan_dep_vld_vec_28[4];
    assign dep_chan_data_28_21 = out_chan_dep_data_28;
    assign token_28_21 = token_out_vec_28[4];
    assign dep_chan_vld_28_22 = out_chan_dep_vld_vec_28[5];
    assign dep_chan_data_28_22 = out_chan_dep_data_28;
    assign token_28_22 = token_out_vec_28[5];
    assign dep_chan_vld_28_23 = out_chan_dep_vld_vec_28[6];
    assign dep_chan_data_28_23 = out_chan_dep_data_28;
    assign token_28_23 = token_out_vec_28[6];
    assign dep_chan_vld_28_24 = out_chan_dep_vld_vec_28[7];
    assign dep_chan_data_28_24 = out_chan_dep_data_28;
    assign token_28_24 = token_out_vec_28[7];
    assign dep_chan_vld_28_25 = out_chan_dep_vld_vec_28[8];
    assign dep_chan_data_28_25 = out_chan_dep_data_28;
    assign token_28_25 = token_out_vec_28[8];
    assign dep_chan_vld_28_26 = out_chan_dep_vld_vec_28[9];
    assign dep_chan_data_28_26 = out_chan_dep_data_28;
    assign token_28_26 = token_out_vec_28[9];
    assign dep_chan_vld_28_27 = out_chan_dep_vld_vec_28[10];
    assign dep_chan_data_28_27 = out_chan_dep_data_28;
    assign token_28_27 = token_out_vec_28[10];
    assign dep_chan_vld_28_29 = out_chan_dep_vld_vec_28[11];
    assign dep_chan_data_28_29 = out_chan_dep_data_28;
    assign token_28_29 = token_out_vec_28[11];
    assign dep_chan_vld_28_30 = out_chan_dep_vld_vec_28[12];
    assign dep_chan_data_28_30 = out_chan_dep_data_28;
    assign token_28_30 = token_out_vec_28[12];
    assign dep_chan_vld_28_31 = out_chan_dep_vld_vec_28[13];
    assign dep_chan_data_28_31 = out_chan_dep_data_28;
    assign token_28_31 = token_out_vec_28[13];
    assign dep_chan_vld_28_32 = out_chan_dep_vld_vec_28[14];
    assign dep_chan_data_28_32 = out_chan_dep_data_28;
    assign token_28_32 = token_out_vec_28[14];
    assign dep_chan_vld_28_33 = out_chan_dep_vld_vec_28[15];
    assign dep_chan_data_28_33 = out_chan_dep_data_28;
    assign token_28_33 = token_out_vec_28[15];
    assign dep_chan_vld_28_34 = out_chan_dep_vld_vec_28[16];
    assign dep_chan_data_28_34 = out_chan_dep_data_28;
    assign token_28_34 = token_out_vec_28[16];

    // Process: write_back58_U0
    kernel_pr_hls_deadlock_detect_unit #(35, 29, 17, 17) kernel_pr_hls_deadlock_detect_unit_29 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_29),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_29),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_29),
        .token_in_vec(token_in_vec_29),
        .dl_detect_in(dl_detect_out),
        .origin(origin[29]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_29),
        .out_chan_dep_data(out_chan_dep_data_29),
        .token_out_vec(token_out_vec_29),
        .dl_detect_out(dl_in_vec[29]));

    assign proc_29_data_FIFO_blk[0] = 1'b0 | (~write_back58_U0.H_blk_n) | (~write_back58_U0.hyperedge_size_blk_n);
    assign proc_29_data_PIPO_blk[0] = 1'b0;
    assign proc_29_start_FIFO_blk[0] = 1'b0 | (~start_for_write_back58_U0_U.if_empty_n & write_back58_U0.ap_idle & ~start_for_write_back58_U0_U.if_write);
    assign proc_29_TLF_FIFO_blk[0] = 1'b0;
    assign proc_29_input_sync_blk[0] = 1'b0;
    assign proc_29_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_29[0] = dl_detect_out ? proc_dep_vld_vec_29_reg[0] : (proc_29_data_FIFO_blk[0] | proc_29_data_PIPO_blk[0] | proc_29_start_FIFO_blk[0] | proc_29_TLF_FIFO_blk[0] | proc_29_input_sync_blk[0] | proc_29_output_sync_blk[0]);
    assign proc_29_data_FIFO_blk[1] = 1'b0 | (~write_back58_U0.value_stream_V_V10_blk_n);
    assign proc_29_data_PIPO_blk[1] = 1'b0;
    assign proc_29_start_FIFO_blk[1] = 1'b0;
    assign proc_29_TLF_FIFO_blk[1] = 1'b0;
    assign proc_29_input_sync_blk[1] = 1'b0;
    assign proc_29_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_29[1] = dl_detect_out ? proc_dep_vld_vec_29_reg[1] : (proc_29_data_FIFO_blk[1] | proc_29_data_PIPO_blk[1] | proc_29_start_FIFO_blk[1] | proc_29_TLF_FIFO_blk[1] | proc_29_input_sync_blk[1] | proc_29_output_sync_blk[1]);
    assign proc_29_data_FIFO_blk[2] = 1'b0;
    assign proc_29_data_PIPO_blk[2] = 1'b0;
    assign proc_29_start_FIFO_blk[2] = 1'b0;
    assign proc_29_TLF_FIFO_blk[2] = 1'b0;
    assign proc_29_input_sync_blk[2] = 1'b0;
    assign proc_29_output_sync_blk[2] = 1'b0 | (ap_done_reg_10 & write_back58_U0.ap_done & ~write_back48_U0.ap_done);
    assign proc_dep_vld_vec_29[2] = dl_detect_out ? proc_dep_vld_vec_29_reg[2] : (proc_29_data_FIFO_blk[2] | proc_29_data_PIPO_blk[2] | proc_29_start_FIFO_blk[2] | proc_29_TLF_FIFO_blk[2] | proc_29_input_sync_blk[2] | proc_29_output_sync_blk[2]);
    assign proc_29_data_FIFO_blk[3] = 1'b0;
    assign proc_29_data_PIPO_blk[3] = 1'b0;
    assign proc_29_start_FIFO_blk[3] = 1'b0;
    assign proc_29_TLF_FIFO_blk[3] = 1'b0;
    assign proc_29_input_sync_blk[3] = 1'b0;
    assign proc_29_output_sync_blk[3] = 1'b0 | (ap_done_reg_10 & write_back58_U0.ap_done & ~write_back49_U0.ap_done);
    assign proc_dep_vld_vec_29[3] = dl_detect_out ? proc_dep_vld_vec_29_reg[3] : (proc_29_data_FIFO_blk[3] | proc_29_data_PIPO_blk[3] | proc_29_start_FIFO_blk[3] | proc_29_TLF_FIFO_blk[3] | proc_29_input_sync_blk[3] | proc_29_output_sync_blk[3]);
    assign proc_29_data_FIFO_blk[4] = 1'b0;
    assign proc_29_data_PIPO_blk[4] = 1'b0;
    assign proc_29_start_FIFO_blk[4] = 1'b0;
    assign proc_29_TLF_FIFO_blk[4] = 1'b0;
    assign proc_29_input_sync_blk[4] = 1'b0;
    assign proc_29_output_sync_blk[4] = 1'b0 | (ap_done_reg_10 & write_back58_U0.ap_done & ~write_back50_U0.ap_done);
    assign proc_dep_vld_vec_29[4] = dl_detect_out ? proc_dep_vld_vec_29_reg[4] : (proc_29_data_FIFO_blk[4] | proc_29_data_PIPO_blk[4] | proc_29_start_FIFO_blk[4] | proc_29_TLF_FIFO_blk[4] | proc_29_input_sync_blk[4] | proc_29_output_sync_blk[4]);
    assign proc_29_data_FIFO_blk[5] = 1'b0;
    assign proc_29_data_PIPO_blk[5] = 1'b0;
    assign proc_29_start_FIFO_blk[5] = 1'b0;
    assign proc_29_TLF_FIFO_blk[5] = 1'b0;
    assign proc_29_input_sync_blk[5] = 1'b0;
    assign proc_29_output_sync_blk[5] = 1'b0 | (ap_done_reg_10 & write_back58_U0.ap_done & ~write_back51_U0.ap_done);
    assign proc_dep_vld_vec_29[5] = dl_detect_out ? proc_dep_vld_vec_29_reg[5] : (proc_29_data_FIFO_blk[5] | proc_29_data_PIPO_blk[5] | proc_29_start_FIFO_blk[5] | proc_29_TLF_FIFO_blk[5] | proc_29_input_sync_blk[5] | proc_29_output_sync_blk[5]);
    assign proc_29_data_FIFO_blk[6] = 1'b0;
    assign proc_29_data_PIPO_blk[6] = 1'b0;
    assign proc_29_start_FIFO_blk[6] = 1'b0;
    assign proc_29_TLF_FIFO_blk[6] = 1'b0;
    assign proc_29_input_sync_blk[6] = 1'b0;
    assign proc_29_output_sync_blk[6] = 1'b0 | (ap_done_reg_10 & write_back58_U0.ap_done & ~write_back52_U0.ap_done);
    assign proc_dep_vld_vec_29[6] = dl_detect_out ? proc_dep_vld_vec_29_reg[6] : (proc_29_data_FIFO_blk[6] | proc_29_data_PIPO_blk[6] | proc_29_start_FIFO_blk[6] | proc_29_TLF_FIFO_blk[6] | proc_29_input_sync_blk[6] | proc_29_output_sync_blk[6]);
    assign proc_29_data_FIFO_blk[7] = 1'b0;
    assign proc_29_data_PIPO_blk[7] = 1'b0;
    assign proc_29_start_FIFO_blk[7] = 1'b0;
    assign proc_29_TLF_FIFO_blk[7] = 1'b0;
    assign proc_29_input_sync_blk[7] = 1'b0;
    assign proc_29_output_sync_blk[7] = 1'b0 | (ap_done_reg_10 & write_back58_U0.ap_done & ~write_back53_U0.ap_done);
    assign proc_dep_vld_vec_29[7] = dl_detect_out ? proc_dep_vld_vec_29_reg[7] : (proc_29_data_FIFO_blk[7] | proc_29_data_PIPO_blk[7] | proc_29_start_FIFO_blk[7] | proc_29_TLF_FIFO_blk[7] | proc_29_input_sync_blk[7] | proc_29_output_sync_blk[7]);
    assign proc_29_data_FIFO_blk[8] = 1'b0;
    assign proc_29_data_PIPO_blk[8] = 1'b0;
    assign proc_29_start_FIFO_blk[8] = 1'b0;
    assign proc_29_TLF_FIFO_blk[8] = 1'b0;
    assign proc_29_input_sync_blk[8] = 1'b0;
    assign proc_29_output_sync_blk[8] = 1'b0 | (ap_done_reg_10 & write_back58_U0.ap_done & ~write_back54_U0.ap_done);
    assign proc_dep_vld_vec_29[8] = dl_detect_out ? proc_dep_vld_vec_29_reg[8] : (proc_29_data_FIFO_blk[8] | proc_29_data_PIPO_blk[8] | proc_29_start_FIFO_blk[8] | proc_29_TLF_FIFO_blk[8] | proc_29_input_sync_blk[8] | proc_29_output_sync_blk[8]);
    assign proc_29_data_FIFO_blk[9] = 1'b0;
    assign proc_29_data_PIPO_blk[9] = 1'b0;
    assign proc_29_start_FIFO_blk[9] = 1'b0;
    assign proc_29_TLF_FIFO_blk[9] = 1'b0;
    assign proc_29_input_sync_blk[9] = 1'b0;
    assign proc_29_output_sync_blk[9] = 1'b0 | (ap_done_reg_10 & write_back58_U0.ap_done & ~write_back55_U0.ap_done);
    assign proc_dep_vld_vec_29[9] = dl_detect_out ? proc_dep_vld_vec_29_reg[9] : (proc_29_data_FIFO_blk[9] | proc_29_data_PIPO_blk[9] | proc_29_start_FIFO_blk[9] | proc_29_TLF_FIFO_blk[9] | proc_29_input_sync_blk[9] | proc_29_output_sync_blk[9]);
    assign proc_29_data_FIFO_blk[10] = 1'b0;
    assign proc_29_data_PIPO_blk[10] = 1'b0;
    assign proc_29_start_FIFO_blk[10] = 1'b0;
    assign proc_29_TLF_FIFO_blk[10] = 1'b0;
    assign proc_29_input_sync_blk[10] = 1'b0;
    assign proc_29_output_sync_blk[10] = 1'b0 | (ap_done_reg_10 & write_back58_U0.ap_done & ~write_back56_U0.ap_done);
    assign proc_dep_vld_vec_29[10] = dl_detect_out ? proc_dep_vld_vec_29_reg[10] : (proc_29_data_FIFO_blk[10] | proc_29_data_PIPO_blk[10] | proc_29_start_FIFO_blk[10] | proc_29_TLF_FIFO_blk[10] | proc_29_input_sync_blk[10] | proc_29_output_sync_blk[10]);
    assign proc_29_data_FIFO_blk[11] = 1'b0;
    assign proc_29_data_PIPO_blk[11] = 1'b0;
    assign proc_29_start_FIFO_blk[11] = 1'b0;
    assign proc_29_TLF_FIFO_blk[11] = 1'b0;
    assign proc_29_input_sync_blk[11] = 1'b0;
    assign proc_29_output_sync_blk[11] = 1'b0 | (ap_done_reg_10 & write_back58_U0.ap_done & ~write_back57_U0.ap_done);
    assign proc_dep_vld_vec_29[11] = dl_detect_out ? proc_dep_vld_vec_29_reg[11] : (proc_29_data_FIFO_blk[11] | proc_29_data_PIPO_blk[11] | proc_29_start_FIFO_blk[11] | proc_29_TLF_FIFO_blk[11] | proc_29_input_sync_blk[11] | proc_29_output_sync_blk[11]);
    assign proc_29_data_FIFO_blk[12] = 1'b0;
    assign proc_29_data_PIPO_blk[12] = 1'b0;
    assign proc_29_start_FIFO_blk[12] = 1'b0;
    assign proc_29_TLF_FIFO_blk[12] = 1'b0;
    assign proc_29_input_sync_blk[12] = 1'b0;
    assign proc_29_output_sync_blk[12] = 1'b0 | (ap_done_reg_10 & write_back58_U0.ap_done & ~write_back59_U0.ap_done);
    assign proc_dep_vld_vec_29[12] = dl_detect_out ? proc_dep_vld_vec_29_reg[12] : (proc_29_data_FIFO_blk[12] | proc_29_data_PIPO_blk[12] | proc_29_start_FIFO_blk[12] | proc_29_TLF_FIFO_blk[12] | proc_29_input_sync_blk[12] | proc_29_output_sync_blk[12]);
    assign proc_29_data_FIFO_blk[13] = 1'b0;
    assign proc_29_data_PIPO_blk[13] = 1'b0;
    assign proc_29_start_FIFO_blk[13] = 1'b0;
    assign proc_29_TLF_FIFO_blk[13] = 1'b0;
    assign proc_29_input_sync_blk[13] = 1'b0;
    assign proc_29_output_sync_blk[13] = 1'b0 | (ap_done_reg_10 & write_back58_U0.ap_done & ~write_back60_U0.ap_done);
    assign proc_dep_vld_vec_29[13] = dl_detect_out ? proc_dep_vld_vec_29_reg[13] : (proc_29_data_FIFO_blk[13] | proc_29_data_PIPO_blk[13] | proc_29_start_FIFO_blk[13] | proc_29_TLF_FIFO_blk[13] | proc_29_input_sync_blk[13] | proc_29_output_sync_blk[13]);
    assign proc_29_data_FIFO_blk[14] = 1'b0;
    assign proc_29_data_PIPO_blk[14] = 1'b0;
    assign proc_29_start_FIFO_blk[14] = 1'b0;
    assign proc_29_TLF_FIFO_blk[14] = 1'b0;
    assign proc_29_input_sync_blk[14] = 1'b0;
    assign proc_29_output_sync_blk[14] = 1'b0 | (ap_done_reg_10 & write_back58_U0.ap_done & ~write_back61_U0.ap_done);
    assign proc_dep_vld_vec_29[14] = dl_detect_out ? proc_dep_vld_vec_29_reg[14] : (proc_29_data_FIFO_blk[14] | proc_29_data_PIPO_blk[14] | proc_29_start_FIFO_blk[14] | proc_29_TLF_FIFO_blk[14] | proc_29_input_sync_blk[14] | proc_29_output_sync_blk[14]);
    assign proc_29_data_FIFO_blk[15] = 1'b0;
    assign proc_29_data_PIPO_blk[15] = 1'b0;
    assign proc_29_start_FIFO_blk[15] = 1'b0;
    assign proc_29_TLF_FIFO_blk[15] = 1'b0;
    assign proc_29_input_sync_blk[15] = 1'b0;
    assign proc_29_output_sync_blk[15] = 1'b0 | (ap_done_reg_10 & write_back58_U0.ap_done & ~write_back62_U0.ap_done);
    assign proc_dep_vld_vec_29[15] = dl_detect_out ? proc_dep_vld_vec_29_reg[15] : (proc_29_data_FIFO_blk[15] | proc_29_data_PIPO_blk[15] | proc_29_start_FIFO_blk[15] | proc_29_TLF_FIFO_blk[15] | proc_29_input_sync_blk[15] | proc_29_output_sync_blk[15]);
    assign proc_29_data_FIFO_blk[16] = 1'b0;
    assign proc_29_data_PIPO_blk[16] = 1'b0;
    assign proc_29_start_FIFO_blk[16] = 1'b0;
    assign proc_29_TLF_FIFO_blk[16] = 1'b0;
    assign proc_29_input_sync_blk[16] = 1'b0;
    assign proc_29_output_sync_blk[16] = 1'b0 | (ap_done_reg_10 & write_back58_U0.ap_done & ~write_back63_U0.ap_done);
    assign proc_dep_vld_vec_29[16] = dl_detect_out ? proc_dep_vld_vec_29_reg[16] : (proc_29_data_FIFO_blk[16] | proc_29_data_PIPO_blk[16] | proc_29_start_FIFO_blk[16] | proc_29_TLF_FIFO_blk[16] | proc_29_input_sync_blk[16] | proc_29_output_sync_blk[16]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_29_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_29_reg <= proc_dep_vld_vec_29;
        end
    end
    assign in_chan_dep_vld_vec_29[0] = dep_chan_vld_0_29;
    assign in_chan_dep_data_vec_29[34 : 0] = dep_chan_data_0_29;
    assign token_in_vec_29[0] = token_0_29;
    assign in_chan_dep_vld_vec_29[1] = dep_chan_vld_13_29;
    assign in_chan_dep_data_vec_29[69 : 35] = dep_chan_data_13_29;
    assign token_in_vec_29[1] = token_13_29;
    assign in_chan_dep_vld_vec_29[2] = dep_chan_vld_19_29;
    assign in_chan_dep_data_vec_29[104 : 70] = dep_chan_data_19_29;
    assign token_in_vec_29[2] = token_19_29;
    assign in_chan_dep_vld_vec_29[3] = dep_chan_vld_20_29;
    assign in_chan_dep_data_vec_29[139 : 105] = dep_chan_data_20_29;
    assign token_in_vec_29[3] = token_20_29;
    assign in_chan_dep_vld_vec_29[4] = dep_chan_vld_21_29;
    assign in_chan_dep_data_vec_29[174 : 140] = dep_chan_data_21_29;
    assign token_in_vec_29[4] = token_21_29;
    assign in_chan_dep_vld_vec_29[5] = dep_chan_vld_22_29;
    assign in_chan_dep_data_vec_29[209 : 175] = dep_chan_data_22_29;
    assign token_in_vec_29[5] = token_22_29;
    assign in_chan_dep_vld_vec_29[6] = dep_chan_vld_23_29;
    assign in_chan_dep_data_vec_29[244 : 210] = dep_chan_data_23_29;
    assign token_in_vec_29[6] = token_23_29;
    assign in_chan_dep_vld_vec_29[7] = dep_chan_vld_24_29;
    assign in_chan_dep_data_vec_29[279 : 245] = dep_chan_data_24_29;
    assign token_in_vec_29[7] = token_24_29;
    assign in_chan_dep_vld_vec_29[8] = dep_chan_vld_25_29;
    assign in_chan_dep_data_vec_29[314 : 280] = dep_chan_data_25_29;
    assign token_in_vec_29[8] = token_25_29;
    assign in_chan_dep_vld_vec_29[9] = dep_chan_vld_26_29;
    assign in_chan_dep_data_vec_29[349 : 315] = dep_chan_data_26_29;
    assign token_in_vec_29[9] = token_26_29;
    assign in_chan_dep_vld_vec_29[10] = dep_chan_vld_27_29;
    assign in_chan_dep_data_vec_29[384 : 350] = dep_chan_data_27_29;
    assign token_in_vec_29[10] = token_27_29;
    assign in_chan_dep_vld_vec_29[11] = dep_chan_vld_28_29;
    assign in_chan_dep_data_vec_29[419 : 385] = dep_chan_data_28_29;
    assign token_in_vec_29[11] = token_28_29;
    assign in_chan_dep_vld_vec_29[12] = dep_chan_vld_30_29;
    assign in_chan_dep_data_vec_29[454 : 420] = dep_chan_data_30_29;
    assign token_in_vec_29[12] = token_30_29;
    assign in_chan_dep_vld_vec_29[13] = dep_chan_vld_31_29;
    assign in_chan_dep_data_vec_29[489 : 455] = dep_chan_data_31_29;
    assign token_in_vec_29[13] = token_31_29;
    assign in_chan_dep_vld_vec_29[14] = dep_chan_vld_32_29;
    assign in_chan_dep_data_vec_29[524 : 490] = dep_chan_data_32_29;
    assign token_in_vec_29[14] = token_32_29;
    assign in_chan_dep_vld_vec_29[15] = dep_chan_vld_33_29;
    assign in_chan_dep_data_vec_29[559 : 525] = dep_chan_data_33_29;
    assign token_in_vec_29[15] = token_33_29;
    assign in_chan_dep_vld_vec_29[16] = dep_chan_vld_34_29;
    assign in_chan_dep_data_vec_29[594 : 560] = dep_chan_data_34_29;
    assign token_in_vec_29[16] = token_34_29;
    assign dep_chan_vld_29_0 = out_chan_dep_vld_vec_29[0];
    assign dep_chan_data_29_0 = out_chan_dep_data_29;
    assign token_29_0 = token_out_vec_29[0];
    assign dep_chan_vld_29_13 = out_chan_dep_vld_vec_29[1];
    assign dep_chan_data_29_13 = out_chan_dep_data_29;
    assign token_29_13 = token_out_vec_29[1];
    assign dep_chan_vld_29_19 = out_chan_dep_vld_vec_29[2];
    assign dep_chan_data_29_19 = out_chan_dep_data_29;
    assign token_29_19 = token_out_vec_29[2];
    assign dep_chan_vld_29_20 = out_chan_dep_vld_vec_29[3];
    assign dep_chan_data_29_20 = out_chan_dep_data_29;
    assign token_29_20 = token_out_vec_29[3];
    assign dep_chan_vld_29_21 = out_chan_dep_vld_vec_29[4];
    assign dep_chan_data_29_21 = out_chan_dep_data_29;
    assign token_29_21 = token_out_vec_29[4];
    assign dep_chan_vld_29_22 = out_chan_dep_vld_vec_29[5];
    assign dep_chan_data_29_22 = out_chan_dep_data_29;
    assign token_29_22 = token_out_vec_29[5];
    assign dep_chan_vld_29_23 = out_chan_dep_vld_vec_29[6];
    assign dep_chan_data_29_23 = out_chan_dep_data_29;
    assign token_29_23 = token_out_vec_29[6];
    assign dep_chan_vld_29_24 = out_chan_dep_vld_vec_29[7];
    assign dep_chan_data_29_24 = out_chan_dep_data_29;
    assign token_29_24 = token_out_vec_29[7];
    assign dep_chan_vld_29_25 = out_chan_dep_vld_vec_29[8];
    assign dep_chan_data_29_25 = out_chan_dep_data_29;
    assign token_29_25 = token_out_vec_29[8];
    assign dep_chan_vld_29_26 = out_chan_dep_vld_vec_29[9];
    assign dep_chan_data_29_26 = out_chan_dep_data_29;
    assign token_29_26 = token_out_vec_29[9];
    assign dep_chan_vld_29_27 = out_chan_dep_vld_vec_29[10];
    assign dep_chan_data_29_27 = out_chan_dep_data_29;
    assign token_29_27 = token_out_vec_29[10];
    assign dep_chan_vld_29_28 = out_chan_dep_vld_vec_29[11];
    assign dep_chan_data_29_28 = out_chan_dep_data_29;
    assign token_29_28 = token_out_vec_29[11];
    assign dep_chan_vld_29_30 = out_chan_dep_vld_vec_29[12];
    assign dep_chan_data_29_30 = out_chan_dep_data_29;
    assign token_29_30 = token_out_vec_29[12];
    assign dep_chan_vld_29_31 = out_chan_dep_vld_vec_29[13];
    assign dep_chan_data_29_31 = out_chan_dep_data_29;
    assign token_29_31 = token_out_vec_29[13];
    assign dep_chan_vld_29_32 = out_chan_dep_vld_vec_29[14];
    assign dep_chan_data_29_32 = out_chan_dep_data_29;
    assign token_29_32 = token_out_vec_29[14];
    assign dep_chan_vld_29_33 = out_chan_dep_vld_vec_29[15];
    assign dep_chan_data_29_33 = out_chan_dep_data_29;
    assign token_29_33 = token_out_vec_29[15];
    assign dep_chan_vld_29_34 = out_chan_dep_vld_vec_29[16];
    assign dep_chan_data_29_34 = out_chan_dep_data_29;
    assign token_29_34 = token_out_vec_29[16];

    // Process: write_back59_U0
    kernel_pr_hls_deadlock_detect_unit #(35, 30, 17, 17) kernel_pr_hls_deadlock_detect_unit_30 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_30),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_30),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_30),
        .token_in_vec(token_in_vec_30),
        .dl_detect_in(dl_detect_out),
        .origin(origin[30]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_30),
        .out_chan_dep_data(out_chan_dep_data_30),
        .token_out_vec(token_out_vec_30),
        .dl_detect_out(dl_in_vec[30]));

    assign proc_30_data_FIFO_blk[0] = 1'b0 | (~write_back59_U0.H_blk_n) | (~write_back59_U0.hyperedge_size_blk_n);
    assign proc_30_data_PIPO_blk[0] = 1'b0;
    assign proc_30_start_FIFO_blk[0] = 1'b0 | (~start_for_write_back59_U0_U.if_empty_n & write_back59_U0.ap_idle & ~start_for_write_back59_U0_U.if_write);
    assign proc_30_TLF_FIFO_blk[0] = 1'b0;
    assign proc_30_input_sync_blk[0] = 1'b0;
    assign proc_30_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_30[0] = dl_detect_out ? proc_dep_vld_vec_30_reg[0] : (proc_30_data_FIFO_blk[0] | proc_30_data_PIPO_blk[0] | proc_30_start_FIFO_blk[0] | proc_30_TLF_FIFO_blk[0] | proc_30_input_sync_blk[0] | proc_30_output_sync_blk[0]);
    assign proc_30_data_FIFO_blk[1] = 1'b0 | (~write_back59_U0.value_stream_V_V11_blk_n);
    assign proc_30_data_PIPO_blk[1] = 1'b0;
    assign proc_30_start_FIFO_blk[1] = 1'b0;
    assign proc_30_TLF_FIFO_blk[1] = 1'b0;
    assign proc_30_input_sync_blk[1] = 1'b0;
    assign proc_30_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_30[1] = dl_detect_out ? proc_dep_vld_vec_30_reg[1] : (proc_30_data_FIFO_blk[1] | proc_30_data_PIPO_blk[1] | proc_30_start_FIFO_blk[1] | proc_30_TLF_FIFO_blk[1] | proc_30_input_sync_blk[1] | proc_30_output_sync_blk[1]);
    assign proc_30_data_FIFO_blk[2] = 1'b0;
    assign proc_30_data_PIPO_blk[2] = 1'b0;
    assign proc_30_start_FIFO_blk[2] = 1'b0;
    assign proc_30_TLF_FIFO_blk[2] = 1'b0;
    assign proc_30_input_sync_blk[2] = 1'b0;
    assign proc_30_output_sync_blk[2] = 1'b0 | (ap_done_reg_11 & write_back59_U0.ap_done & ~write_back48_U0.ap_done);
    assign proc_dep_vld_vec_30[2] = dl_detect_out ? proc_dep_vld_vec_30_reg[2] : (proc_30_data_FIFO_blk[2] | proc_30_data_PIPO_blk[2] | proc_30_start_FIFO_blk[2] | proc_30_TLF_FIFO_blk[2] | proc_30_input_sync_blk[2] | proc_30_output_sync_blk[2]);
    assign proc_30_data_FIFO_blk[3] = 1'b0;
    assign proc_30_data_PIPO_blk[3] = 1'b0;
    assign proc_30_start_FIFO_blk[3] = 1'b0;
    assign proc_30_TLF_FIFO_blk[3] = 1'b0;
    assign proc_30_input_sync_blk[3] = 1'b0;
    assign proc_30_output_sync_blk[3] = 1'b0 | (ap_done_reg_11 & write_back59_U0.ap_done & ~write_back49_U0.ap_done);
    assign proc_dep_vld_vec_30[3] = dl_detect_out ? proc_dep_vld_vec_30_reg[3] : (proc_30_data_FIFO_blk[3] | proc_30_data_PIPO_blk[3] | proc_30_start_FIFO_blk[3] | proc_30_TLF_FIFO_blk[3] | proc_30_input_sync_blk[3] | proc_30_output_sync_blk[3]);
    assign proc_30_data_FIFO_blk[4] = 1'b0;
    assign proc_30_data_PIPO_blk[4] = 1'b0;
    assign proc_30_start_FIFO_blk[4] = 1'b0;
    assign proc_30_TLF_FIFO_blk[4] = 1'b0;
    assign proc_30_input_sync_blk[4] = 1'b0;
    assign proc_30_output_sync_blk[4] = 1'b0 | (ap_done_reg_11 & write_back59_U0.ap_done & ~write_back50_U0.ap_done);
    assign proc_dep_vld_vec_30[4] = dl_detect_out ? proc_dep_vld_vec_30_reg[4] : (proc_30_data_FIFO_blk[4] | proc_30_data_PIPO_blk[4] | proc_30_start_FIFO_blk[4] | proc_30_TLF_FIFO_blk[4] | proc_30_input_sync_blk[4] | proc_30_output_sync_blk[4]);
    assign proc_30_data_FIFO_blk[5] = 1'b0;
    assign proc_30_data_PIPO_blk[5] = 1'b0;
    assign proc_30_start_FIFO_blk[5] = 1'b0;
    assign proc_30_TLF_FIFO_blk[5] = 1'b0;
    assign proc_30_input_sync_blk[5] = 1'b0;
    assign proc_30_output_sync_blk[5] = 1'b0 | (ap_done_reg_11 & write_back59_U0.ap_done & ~write_back51_U0.ap_done);
    assign proc_dep_vld_vec_30[5] = dl_detect_out ? proc_dep_vld_vec_30_reg[5] : (proc_30_data_FIFO_blk[5] | proc_30_data_PIPO_blk[5] | proc_30_start_FIFO_blk[5] | proc_30_TLF_FIFO_blk[5] | proc_30_input_sync_blk[5] | proc_30_output_sync_blk[5]);
    assign proc_30_data_FIFO_blk[6] = 1'b0;
    assign proc_30_data_PIPO_blk[6] = 1'b0;
    assign proc_30_start_FIFO_blk[6] = 1'b0;
    assign proc_30_TLF_FIFO_blk[6] = 1'b0;
    assign proc_30_input_sync_blk[6] = 1'b0;
    assign proc_30_output_sync_blk[6] = 1'b0 | (ap_done_reg_11 & write_back59_U0.ap_done & ~write_back52_U0.ap_done);
    assign proc_dep_vld_vec_30[6] = dl_detect_out ? proc_dep_vld_vec_30_reg[6] : (proc_30_data_FIFO_blk[6] | proc_30_data_PIPO_blk[6] | proc_30_start_FIFO_blk[6] | proc_30_TLF_FIFO_blk[6] | proc_30_input_sync_blk[6] | proc_30_output_sync_blk[6]);
    assign proc_30_data_FIFO_blk[7] = 1'b0;
    assign proc_30_data_PIPO_blk[7] = 1'b0;
    assign proc_30_start_FIFO_blk[7] = 1'b0;
    assign proc_30_TLF_FIFO_blk[7] = 1'b0;
    assign proc_30_input_sync_blk[7] = 1'b0;
    assign proc_30_output_sync_blk[7] = 1'b0 | (ap_done_reg_11 & write_back59_U0.ap_done & ~write_back53_U0.ap_done);
    assign proc_dep_vld_vec_30[7] = dl_detect_out ? proc_dep_vld_vec_30_reg[7] : (proc_30_data_FIFO_blk[7] | proc_30_data_PIPO_blk[7] | proc_30_start_FIFO_blk[7] | proc_30_TLF_FIFO_blk[7] | proc_30_input_sync_blk[7] | proc_30_output_sync_blk[7]);
    assign proc_30_data_FIFO_blk[8] = 1'b0;
    assign proc_30_data_PIPO_blk[8] = 1'b0;
    assign proc_30_start_FIFO_blk[8] = 1'b0;
    assign proc_30_TLF_FIFO_blk[8] = 1'b0;
    assign proc_30_input_sync_blk[8] = 1'b0;
    assign proc_30_output_sync_blk[8] = 1'b0 | (ap_done_reg_11 & write_back59_U0.ap_done & ~write_back54_U0.ap_done);
    assign proc_dep_vld_vec_30[8] = dl_detect_out ? proc_dep_vld_vec_30_reg[8] : (proc_30_data_FIFO_blk[8] | proc_30_data_PIPO_blk[8] | proc_30_start_FIFO_blk[8] | proc_30_TLF_FIFO_blk[8] | proc_30_input_sync_blk[8] | proc_30_output_sync_blk[8]);
    assign proc_30_data_FIFO_blk[9] = 1'b0;
    assign proc_30_data_PIPO_blk[9] = 1'b0;
    assign proc_30_start_FIFO_blk[9] = 1'b0;
    assign proc_30_TLF_FIFO_blk[9] = 1'b0;
    assign proc_30_input_sync_blk[9] = 1'b0;
    assign proc_30_output_sync_blk[9] = 1'b0 | (ap_done_reg_11 & write_back59_U0.ap_done & ~write_back55_U0.ap_done);
    assign proc_dep_vld_vec_30[9] = dl_detect_out ? proc_dep_vld_vec_30_reg[9] : (proc_30_data_FIFO_blk[9] | proc_30_data_PIPO_blk[9] | proc_30_start_FIFO_blk[9] | proc_30_TLF_FIFO_blk[9] | proc_30_input_sync_blk[9] | proc_30_output_sync_blk[9]);
    assign proc_30_data_FIFO_blk[10] = 1'b0;
    assign proc_30_data_PIPO_blk[10] = 1'b0;
    assign proc_30_start_FIFO_blk[10] = 1'b0;
    assign proc_30_TLF_FIFO_blk[10] = 1'b0;
    assign proc_30_input_sync_blk[10] = 1'b0;
    assign proc_30_output_sync_blk[10] = 1'b0 | (ap_done_reg_11 & write_back59_U0.ap_done & ~write_back56_U0.ap_done);
    assign proc_dep_vld_vec_30[10] = dl_detect_out ? proc_dep_vld_vec_30_reg[10] : (proc_30_data_FIFO_blk[10] | proc_30_data_PIPO_blk[10] | proc_30_start_FIFO_blk[10] | proc_30_TLF_FIFO_blk[10] | proc_30_input_sync_blk[10] | proc_30_output_sync_blk[10]);
    assign proc_30_data_FIFO_blk[11] = 1'b0;
    assign proc_30_data_PIPO_blk[11] = 1'b0;
    assign proc_30_start_FIFO_blk[11] = 1'b0;
    assign proc_30_TLF_FIFO_blk[11] = 1'b0;
    assign proc_30_input_sync_blk[11] = 1'b0;
    assign proc_30_output_sync_blk[11] = 1'b0 | (ap_done_reg_11 & write_back59_U0.ap_done & ~write_back57_U0.ap_done);
    assign proc_dep_vld_vec_30[11] = dl_detect_out ? proc_dep_vld_vec_30_reg[11] : (proc_30_data_FIFO_blk[11] | proc_30_data_PIPO_blk[11] | proc_30_start_FIFO_blk[11] | proc_30_TLF_FIFO_blk[11] | proc_30_input_sync_blk[11] | proc_30_output_sync_blk[11]);
    assign proc_30_data_FIFO_blk[12] = 1'b0;
    assign proc_30_data_PIPO_blk[12] = 1'b0;
    assign proc_30_start_FIFO_blk[12] = 1'b0;
    assign proc_30_TLF_FIFO_blk[12] = 1'b0;
    assign proc_30_input_sync_blk[12] = 1'b0;
    assign proc_30_output_sync_blk[12] = 1'b0 | (ap_done_reg_11 & write_back59_U0.ap_done & ~write_back58_U0.ap_done);
    assign proc_dep_vld_vec_30[12] = dl_detect_out ? proc_dep_vld_vec_30_reg[12] : (proc_30_data_FIFO_blk[12] | proc_30_data_PIPO_blk[12] | proc_30_start_FIFO_blk[12] | proc_30_TLF_FIFO_blk[12] | proc_30_input_sync_blk[12] | proc_30_output_sync_blk[12]);
    assign proc_30_data_FIFO_blk[13] = 1'b0;
    assign proc_30_data_PIPO_blk[13] = 1'b0;
    assign proc_30_start_FIFO_blk[13] = 1'b0;
    assign proc_30_TLF_FIFO_blk[13] = 1'b0;
    assign proc_30_input_sync_blk[13] = 1'b0;
    assign proc_30_output_sync_blk[13] = 1'b0 | (ap_done_reg_11 & write_back59_U0.ap_done & ~write_back60_U0.ap_done);
    assign proc_dep_vld_vec_30[13] = dl_detect_out ? proc_dep_vld_vec_30_reg[13] : (proc_30_data_FIFO_blk[13] | proc_30_data_PIPO_blk[13] | proc_30_start_FIFO_blk[13] | proc_30_TLF_FIFO_blk[13] | proc_30_input_sync_blk[13] | proc_30_output_sync_blk[13]);
    assign proc_30_data_FIFO_blk[14] = 1'b0;
    assign proc_30_data_PIPO_blk[14] = 1'b0;
    assign proc_30_start_FIFO_blk[14] = 1'b0;
    assign proc_30_TLF_FIFO_blk[14] = 1'b0;
    assign proc_30_input_sync_blk[14] = 1'b0;
    assign proc_30_output_sync_blk[14] = 1'b0 | (ap_done_reg_11 & write_back59_U0.ap_done & ~write_back61_U0.ap_done);
    assign proc_dep_vld_vec_30[14] = dl_detect_out ? proc_dep_vld_vec_30_reg[14] : (proc_30_data_FIFO_blk[14] | proc_30_data_PIPO_blk[14] | proc_30_start_FIFO_blk[14] | proc_30_TLF_FIFO_blk[14] | proc_30_input_sync_blk[14] | proc_30_output_sync_blk[14]);
    assign proc_30_data_FIFO_blk[15] = 1'b0;
    assign proc_30_data_PIPO_blk[15] = 1'b0;
    assign proc_30_start_FIFO_blk[15] = 1'b0;
    assign proc_30_TLF_FIFO_blk[15] = 1'b0;
    assign proc_30_input_sync_blk[15] = 1'b0;
    assign proc_30_output_sync_blk[15] = 1'b0 | (ap_done_reg_11 & write_back59_U0.ap_done & ~write_back62_U0.ap_done);
    assign proc_dep_vld_vec_30[15] = dl_detect_out ? proc_dep_vld_vec_30_reg[15] : (proc_30_data_FIFO_blk[15] | proc_30_data_PIPO_blk[15] | proc_30_start_FIFO_blk[15] | proc_30_TLF_FIFO_blk[15] | proc_30_input_sync_blk[15] | proc_30_output_sync_blk[15]);
    assign proc_30_data_FIFO_blk[16] = 1'b0;
    assign proc_30_data_PIPO_blk[16] = 1'b0;
    assign proc_30_start_FIFO_blk[16] = 1'b0;
    assign proc_30_TLF_FIFO_blk[16] = 1'b0;
    assign proc_30_input_sync_blk[16] = 1'b0;
    assign proc_30_output_sync_blk[16] = 1'b0 | (ap_done_reg_11 & write_back59_U0.ap_done & ~write_back63_U0.ap_done);
    assign proc_dep_vld_vec_30[16] = dl_detect_out ? proc_dep_vld_vec_30_reg[16] : (proc_30_data_FIFO_blk[16] | proc_30_data_PIPO_blk[16] | proc_30_start_FIFO_blk[16] | proc_30_TLF_FIFO_blk[16] | proc_30_input_sync_blk[16] | proc_30_output_sync_blk[16]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_30_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_30_reg <= proc_dep_vld_vec_30;
        end
    end
    assign in_chan_dep_vld_vec_30[0] = dep_chan_vld_0_30;
    assign in_chan_dep_data_vec_30[34 : 0] = dep_chan_data_0_30;
    assign token_in_vec_30[0] = token_0_30;
    assign in_chan_dep_vld_vec_30[1] = dep_chan_vld_14_30;
    assign in_chan_dep_data_vec_30[69 : 35] = dep_chan_data_14_30;
    assign token_in_vec_30[1] = token_14_30;
    assign in_chan_dep_vld_vec_30[2] = dep_chan_vld_19_30;
    assign in_chan_dep_data_vec_30[104 : 70] = dep_chan_data_19_30;
    assign token_in_vec_30[2] = token_19_30;
    assign in_chan_dep_vld_vec_30[3] = dep_chan_vld_20_30;
    assign in_chan_dep_data_vec_30[139 : 105] = dep_chan_data_20_30;
    assign token_in_vec_30[3] = token_20_30;
    assign in_chan_dep_vld_vec_30[4] = dep_chan_vld_21_30;
    assign in_chan_dep_data_vec_30[174 : 140] = dep_chan_data_21_30;
    assign token_in_vec_30[4] = token_21_30;
    assign in_chan_dep_vld_vec_30[5] = dep_chan_vld_22_30;
    assign in_chan_dep_data_vec_30[209 : 175] = dep_chan_data_22_30;
    assign token_in_vec_30[5] = token_22_30;
    assign in_chan_dep_vld_vec_30[6] = dep_chan_vld_23_30;
    assign in_chan_dep_data_vec_30[244 : 210] = dep_chan_data_23_30;
    assign token_in_vec_30[6] = token_23_30;
    assign in_chan_dep_vld_vec_30[7] = dep_chan_vld_24_30;
    assign in_chan_dep_data_vec_30[279 : 245] = dep_chan_data_24_30;
    assign token_in_vec_30[7] = token_24_30;
    assign in_chan_dep_vld_vec_30[8] = dep_chan_vld_25_30;
    assign in_chan_dep_data_vec_30[314 : 280] = dep_chan_data_25_30;
    assign token_in_vec_30[8] = token_25_30;
    assign in_chan_dep_vld_vec_30[9] = dep_chan_vld_26_30;
    assign in_chan_dep_data_vec_30[349 : 315] = dep_chan_data_26_30;
    assign token_in_vec_30[9] = token_26_30;
    assign in_chan_dep_vld_vec_30[10] = dep_chan_vld_27_30;
    assign in_chan_dep_data_vec_30[384 : 350] = dep_chan_data_27_30;
    assign token_in_vec_30[10] = token_27_30;
    assign in_chan_dep_vld_vec_30[11] = dep_chan_vld_28_30;
    assign in_chan_dep_data_vec_30[419 : 385] = dep_chan_data_28_30;
    assign token_in_vec_30[11] = token_28_30;
    assign in_chan_dep_vld_vec_30[12] = dep_chan_vld_29_30;
    assign in_chan_dep_data_vec_30[454 : 420] = dep_chan_data_29_30;
    assign token_in_vec_30[12] = token_29_30;
    assign in_chan_dep_vld_vec_30[13] = dep_chan_vld_31_30;
    assign in_chan_dep_data_vec_30[489 : 455] = dep_chan_data_31_30;
    assign token_in_vec_30[13] = token_31_30;
    assign in_chan_dep_vld_vec_30[14] = dep_chan_vld_32_30;
    assign in_chan_dep_data_vec_30[524 : 490] = dep_chan_data_32_30;
    assign token_in_vec_30[14] = token_32_30;
    assign in_chan_dep_vld_vec_30[15] = dep_chan_vld_33_30;
    assign in_chan_dep_data_vec_30[559 : 525] = dep_chan_data_33_30;
    assign token_in_vec_30[15] = token_33_30;
    assign in_chan_dep_vld_vec_30[16] = dep_chan_vld_34_30;
    assign in_chan_dep_data_vec_30[594 : 560] = dep_chan_data_34_30;
    assign token_in_vec_30[16] = token_34_30;
    assign dep_chan_vld_30_0 = out_chan_dep_vld_vec_30[0];
    assign dep_chan_data_30_0 = out_chan_dep_data_30;
    assign token_30_0 = token_out_vec_30[0];
    assign dep_chan_vld_30_14 = out_chan_dep_vld_vec_30[1];
    assign dep_chan_data_30_14 = out_chan_dep_data_30;
    assign token_30_14 = token_out_vec_30[1];
    assign dep_chan_vld_30_19 = out_chan_dep_vld_vec_30[2];
    assign dep_chan_data_30_19 = out_chan_dep_data_30;
    assign token_30_19 = token_out_vec_30[2];
    assign dep_chan_vld_30_20 = out_chan_dep_vld_vec_30[3];
    assign dep_chan_data_30_20 = out_chan_dep_data_30;
    assign token_30_20 = token_out_vec_30[3];
    assign dep_chan_vld_30_21 = out_chan_dep_vld_vec_30[4];
    assign dep_chan_data_30_21 = out_chan_dep_data_30;
    assign token_30_21 = token_out_vec_30[4];
    assign dep_chan_vld_30_22 = out_chan_dep_vld_vec_30[5];
    assign dep_chan_data_30_22 = out_chan_dep_data_30;
    assign token_30_22 = token_out_vec_30[5];
    assign dep_chan_vld_30_23 = out_chan_dep_vld_vec_30[6];
    assign dep_chan_data_30_23 = out_chan_dep_data_30;
    assign token_30_23 = token_out_vec_30[6];
    assign dep_chan_vld_30_24 = out_chan_dep_vld_vec_30[7];
    assign dep_chan_data_30_24 = out_chan_dep_data_30;
    assign token_30_24 = token_out_vec_30[7];
    assign dep_chan_vld_30_25 = out_chan_dep_vld_vec_30[8];
    assign dep_chan_data_30_25 = out_chan_dep_data_30;
    assign token_30_25 = token_out_vec_30[8];
    assign dep_chan_vld_30_26 = out_chan_dep_vld_vec_30[9];
    assign dep_chan_data_30_26 = out_chan_dep_data_30;
    assign token_30_26 = token_out_vec_30[9];
    assign dep_chan_vld_30_27 = out_chan_dep_vld_vec_30[10];
    assign dep_chan_data_30_27 = out_chan_dep_data_30;
    assign token_30_27 = token_out_vec_30[10];
    assign dep_chan_vld_30_28 = out_chan_dep_vld_vec_30[11];
    assign dep_chan_data_30_28 = out_chan_dep_data_30;
    assign token_30_28 = token_out_vec_30[11];
    assign dep_chan_vld_30_29 = out_chan_dep_vld_vec_30[12];
    assign dep_chan_data_30_29 = out_chan_dep_data_30;
    assign token_30_29 = token_out_vec_30[12];
    assign dep_chan_vld_30_31 = out_chan_dep_vld_vec_30[13];
    assign dep_chan_data_30_31 = out_chan_dep_data_30;
    assign token_30_31 = token_out_vec_30[13];
    assign dep_chan_vld_30_32 = out_chan_dep_vld_vec_30[14];
    assign dep_chan_data_30_32 = out_chan_dep_data_30;
    assign token_30_32 = token_out_vec_30[14];
    assign dep_chan_vld_30_33 = out_chan_dep_vld_vec_30[15];
    assign dep_chan_data_30_33 = out_chan_dep_data_30;
    assign token_30_33 = token_out_vec_30[15];
    assign dep_chan_vld_30_34 = out_chan_dep_vld_vec_30[16];
    assign dep_chan_data_30_34 = out_chan_dep_data_30;
    assign token_30_34 = token_out_vec_30[16];

    // Process: write_back60_U0
    kernel_pr_hls_deadlock_detect_unit #(35, 31, 17, 17) kernel_pr_hls_deadlock_detect_unit_31 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_31),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_31),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_31),
        .token_in_vec(token_in_vec_31),
        .dl_detect_in(dl_detect_out),
        .origin(origin[31]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_31),
        .out_chan_dep_data(out_chan_dep_data_31),
        .token_out_vec(token_out_vec_31),
        .dl_detect_out(dl_in_vec[31]));

    assign proc_31_data_FIFO_blk[0] = 1'b0 | (~write_back60_U0.H_blk_n) | (~write_back60_U0.hyperedge_size_blk_n);
    assign proc_31_data_PIPO_blk[0] = 1'b0;
    assign proc_31_start_FIFO_blk[0] = 1'b0 | (~start_for_write_back60_U0_U.if_empty_n & write_back60_U0.ap_idle & ~start_for_write_back60_U0_U.if_write);
    assign proc_31_TLF_FIFO_blk[0] = 1'b0;
    assign proc_31_input_sync_blk[0] = 1'b0;
    assign proc_31_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_31[0] = dl_detect_out ? proc_dep_vld_vec_31_reg[0] : (proc_31_data_FIFO_blk[0] | proc_31_data_PIPO_blk[0] | proc_31_start_FIFO_blk[0] | proc_31_TLF_FIFO_blk[0] | proc_31_input_sync_blk[0] | proc_31_output_sync_blk[0]);
    assign proc_31_data_FIFO_blk[1] = 1'b0 | (~write_back60_U0.value_stream_V_V12_blk_n);
    assign proc_31_data_PIPO_blk[1] = 1'b0;
    assign proc_31_start_FIFO_blk[1] = 1'b0;
    assign proc_31_TLF_FIFO_blk[1] = 1'b0;
    assign proc_31_input_sync_blk[1] = 1'b0;
    assign proc_31_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_31[1] = dl_detect_out ? proc_dep_vld_vec_31_reg[1] : (proc_31_data_FIFO_blk[1] | proc_31_data_PIPO_blk[1] | proc_31_start_FIFO_blk[1] | proc_31_TLF_FIFO_blk[1] | proc_31_input_sync_blk[1] | proc_31_output_sync_blk[1]);
    assign proc_31_data_FIFO_blk[2] = 1'b0;
    assign proc_31_data_PIPO_blk[2] = 1'b0;
    assign proc_31_start_FIFO_blk[2] = 1'b0;
    assign proc_31_TLF_FIFO_blk[2] = 1'b0;
    assign proc_31_input_sync_blk[2] = 1'b0;
    assign proc_31_output_sync_blk[2] = 1'b0 | (ap_done_reg_12 & write_back60_U0.ap_done & ~write_back48_U0.ap_done);
    assign proc_dep_vld_vec_31[2] = dl_detect_out ? proc_dep_vld_vec_31_reg[2] : (proc_31_data_FIFO_blk[2] | proc_31_data_PIPO_blk[2] | proc_31_start_FIFO_blk[2] | proc_31_TLF_FIFO_blk[2] | proc_31_input_sync_blk[2] | proc_31_output_sync_blk[2]);
    assign proc_31_data_FIFO_blk[3] = 1'b0;
    assign proc_31_data_PIPO_blk[3] = 1'b0;
    assign proc_31_start_FIFO_blk[3] = 1'b0;
    assign proc_31_TLF_FIFO_blk[3] = 1'b0;
    assign proc_31_input_sync_blk[3] = 1'b0;
    assign proc_31_output_sync_blk[3] = 1'b0 | (ap_done_reg_12 & write_back60_U0.ap_done & ~write_back49_U0.ap_done);
    assign proc_dep_vld_vec_31[3] = dl_detect_out ? proc_dep_vld_vec_31_reg[3] : (proc_31_data_FIFO_blk[3] | proc_31_data_PIPO_blk[3] | proc_31_start_FIFO_blk[3] | proc_31_TLF_FIFO_blk[3] | proc_31_input_sync_blk[3] | proc_31_output_sync_blk[3]);
    assign proc_31_data_FIFO_blk[4] = 1'b0;
    assign proc_31_data_PIPO_blk[4] = 1'b0;
    assign proc_31_start_FIFO_blk[4] = 1'b0;
    assign proc_31_TLF_FIFO_blk[4] = 1'b0;
    assign proc_31_input_sync_blk[4] = 1'b0;
    assign proc_31_output_sync_blk[4] = 1'b0 | (ap_done_reg_12 & write_back60_U0.ap_done & ~write_back50_U0.ap_done);
    assign proc_dep_vld_vec_31[4] = dl_detect_out ? proc_dep_vld_vec_31_reg[4] : (proc_31_data_FIFO_blk[4] | proc_31_data_PIPO_blk[4] | proc_31_start_FIFO_blk[4] | proc_31_TLF_FIFO_blk[4] | proc_31_input_sync_blk[4] | proc_31_output_sync_blk[4]);
    assign proc_31_data_FIFO_blk[5] = 1'b0;
    assign proc_31_data_PIPO_blk[5] = 1'b0;
    assign proc_31_start_FIFO_blk[5] = 1'b0;
    assign proc_31_TLF_FIFO_blk[5] = 1'b0;
    assign proc_31_input_sync_blk[5] = 1'b0;
    assign proc_31_output_sync_blk[5] = 1'b0 | (ap_done_reg_12 & write_back60_U0.ap_done & ~write_back51_U0.ap_done);
    assign proc_dep_vld_vec_31[5] = dl_detect_out ? proc_dep_vld_vec_31_reg[5] : (proc_31_data_FIFO_blk[5] | proc_31_data_PIPO_blk[5] | proc_31_start_FIFO_blk[5] | proc_31_TLF_FIFO_blk[5] | proc_31_input_sync_blk[5] | proc_31_output_sync_blk[5]);
    assign proc_31_data_FIFO_blk[6] = 1'b0;
    assign proc_31_data_PIPO_blk[6] = 1'b0;
    assign proc_31_start_FIFO_blk[6] = 1'b0;
    assign proc_31_TLF_FIFO_blk[6] = 1'b0;
    assign proc_31_input_sync_blk[6] = 1'b0;
    assign proc_31_output_sync_blk[6] = 1'b0 | (ap_done_reg_12 & write_back60_U0.ap_done & ~write_back52_U0.ap_done);
    assign proc_dep_vld_vec_31[6] = dl_detect_out ? proc_dep_vld_vec_31_reg[6] : (proc_31_data_FIFO_blk[6] | proc_31_data_PIPO_blk[6] | proc_31_start_FIFO_blk[6] | proc_31_TLF_FIFO_blk[6] | proc_31_input_sync_blk[6] | proc_31_output_sync_blk[6]);
    assign proc_31_data_FIFO_blk[7] = 1'b0;
    assign proc_31_data_PIPO_blk[7] = 1'b0;
    assign proc_31_start_FIFO_blk[7] = 1'b0;
    assign proc_31_TLF_FIFO_blk[7] = 1'b0;
    assign proc_31_input_sync_blk[7] = 1'b0;
    assign proc_31_output_sync_blk[7] = 1'b0 | (ap_done_reg_12 & write_back60_U0.ap_done & ~write_back53_U0.ap_done);
    assign proc_dep_vld_vec_31[7] = dl_detect_out ? proc_dep_vld_vec_31_reg[7] : (proc_31_data_FIFO_blk[7] | proc_31_data_PIPO_blk[7] | proc_31_start_FIFO_blk[7] | proc_31_TLF_FIFO_blk[7] | proc_31_input_sync_blk[7] | proc_31_output_sync_blk[7]);
    assign proc_31_data_FIFO_blk[8] = 1'b0;
    assign proc_31_data_PIPO_blk[8] = 1'b0;
    assign proc_31_start_FIFO_blk[8] = 1'b0;
    assign proc_31_TLF_FIFO_blk[8] = 1'b0;
    assign proc_31_input_sync_blk[8] = 1'b0;
    assign proc_31_output_sync_blk[8] = 1'b0 | (ap_done_reg_12 & write_back60_U0.ap_done & ~write_back54_U0.ap_done);
    assign proc_dep_vld_vec_31[8] = dl_detect_out ? proc_dep_vld_vec_31_reg[8] : (proc_31_data_FIFO_blk[8] | proc_31_data_PIPO_blk[8] | proc_31_start_FIFO_blk[8] | proc_31_TLF_FIFO_blk[8] | proc_31_input_sync_blk[8] | proc_31_output_sync_blk[8]);
    assign proc_31_data_FIFO_blk[9] = 1'b0;
    assign proc_31_data_PIPO_blk[9] = 1'b0;
    assign proc_31_start_FIFO_blk[9] = 1'b0;
    assign proc_31_TLF_FIFO_blk[9] = 1'b0;
    assign proc_31_input_sync_blk[9] = 1'b0;
    assign proc_31_output_sync_blk[9] = 1'b0 | (ap_done_reg_12 & write_back60_U0.ap_done & ~write_back55_U0.ap_done);
    assign proc_dep_vld_vec_31[9] = dl_detect_out ? proc_dep_vld_vec_31_reg[9] : (proc_31_data_FIFO_blk[9] | proc_31_data_PIPO_blk[9] | proc_31_start_FIFO_blk[9] | proc_31_TLF_FIFO_blk[9] | proc_31_input_sync_blk[9] | proc_31_output_sync_blk[9]);
    assign proc_31_data_FIFO_blk[10] = 1'b0;
    assign proc_31_data_PIPO_blk[10] = 1'b0;
    assign proc_31_start_FIFO_blk[10] = 1'b0;
    assign proc_31_TLF_FIFO_blk[10] = 1'b0;
    assign proc_31_input_sync_blk[10] = 1'b0;
    assign proc_31_output_sync_blk[10] = 1'b0 | (ap_done_reg_12 & write_back60_U0.ap_done & ~write_back56_U0.ap_done);
    assign proc_dep_vld_vec_31[10] = dl_detect_out ? proc_dep_vld_vec_31_reg[10] : (proc_31_data_FIFO_blk[10] | proc_31_data_PIPO_blk[10] | proc_31_start_FIFO_blk[10] | proc_31_TLF_FIFO_blk[10] | proc_31_input_sync_blk[10] | proc_31_output_sync_blk[10]);
    assign proc_31_data_FIFO_blk[11] = 1'b0;
    assign proc_31_data_PIPO_blk[11] = 1'b0;
    assign proc_31_start_FIFO_blk[11] = 1'b0;
    assign proc_31_TLF_FIFO_blk[11] = 1'b0;
    assign proc_31_input_sync_blk[11] = 1'b0;
    assign proc_31_output_sync_blk[11] = 1'b0 | (ap_done_reg_12 & write_back60_U0.ap_done & ~write_back57_U0.ap_done);
    assign proc_dep_vld_vec_31[11] = dl_detect_out ? proc_dep_vld_vec_31_reg[11] : (proc_31_data_FIFO_blk[11] | proc_31_data_PIPO_blk[11] | proc_31_start_FIFO_blk[11] | proc_31_TLF_FIFO_blk[11] | proc_31_input_sync_blk[11] | proc_31_output_sync_blk[11]);
    assign proc_31_data_FIFO_blk[12] = 1'b0;
    assign proc_31_data_PIPO_blk[12] = 1'b0;
    assign proc_31_start_FIFO_blk[12] = 1'b0;
    assign proc_31_TLF_FIFO_blk[12] = 1'b0;
    assign proc_31_input_sync_blk[12] = 1'b0;
    assign proc_31_output_sync_blk[12] = 1'b0 | (ap_done_reg_12 & write_back60_U0.ap_done & ~write_back58_U0.ap_done);
    assign proc_dep_vld_vec_31[12] = dl_detect_out ? proc_dep_vld_vec_31_reg[12] : (proc_31_data_FIFO_blk[12] | proc_31_data_PIPO_blk[12] | proc_31_start_FIFO_blk[12] | proc_31_TLF_FIFO_blk[12] | proc_31_input_sync_blk[12] | proc_31_output_sync_blk[12]);
    assign proc_31_data_FIFO_blk[13] = 1'b0;
    assign proc_31_data_PIPO_blk[13] = 1'b0;
    assign proc_31_start_FIFO_blk[13] = 1'b0;
    assign proc_31_TLF_FIFO_blk[13] = 1'b0;
    assign proc_31_input_sync_blk[13] = 1'b0;
    assign proc_31_output_sync_blk[13] = 1'b0 | (ap_done_reg_12 & write_back60_U0.ap_done & ~write_back59_U0.ap_done);
    assign proc_dep_vld_vec_31[13] = dl_detect_out ? proc_dep_vld_vec_31_reg[13] : (proc_31_data_FIFO_blk[13] | proc_31_data_PIPO_blk[13] | proc_31_start_FIFO_blk[13] | proc_31_TLF_FIFO_blk[13] | proc_31_input_sync_blk[13] | proc_31_output_sync_blk[13]);
    assign proc_31_data_FIFO_blk[14] = 1'b0;
    assign proc_31_data_PIPO_blk[14] = 1'b0;
    assign proc_31_start_FIFO_blk[14] = 1'b0;
    assign proc_31_TLF_FIFO_blk[14] = 1'b0;
    assign proc_31_input_sync_blk[14] = 1'b0;
    assign proc_31_output_sync_blk[14] = 1'b0 | (ap_done_reg_12 & write_back60_U0.ap_done & ~write_back61_U0.ap_done);
    assign proc_dep_vld_vec_31[14] = dl_detect_out ? proc_dep_vld_vec_31_reg[14] : (proc_31_data_FIFO_blk[14] | proc_31_data_PIPO_blk[14] | proc_31_start_FIFO_blk[14] | proc_31_TLF_FIFO_blk[14] | proc_31_input_sync_blk[14] | proc_31_output_sync_blk[14]);
    assign proc_31_data_FIFO_blk[15] = 1'b0;
    assign proc_31_data_PIPO_blk[15] = 1'b0;
    assign proc_31_start_FIFO_blk[15] = 1'b0;
    assign proc_31_TLF_FIFO_blk[15] = 1'b0;
    assign proc_31_input_sync_blk[15] = 1'b0;
    assign proc_31_output_sync_blk[15] = 1'b0 | (ap_done_reg_12 & write_back60_U0.ap_done & ~write_back62_U0.ap_done);
    assign proc_dep_vld_vec_31[15] = dl_detect_out ? proc_dep_vld_vec_31_reg[15] : (proc_31_data_FIFO_blk[15] | proc_31_data_PIPO_blk[15] | proc_31_start_FIFO_blk[15] | proc_31_TLF_FIFO_blk[15] | proc_31_input_sync_blk[15] | proc_31_output_sync_blk[15]);
    assign proc_31_data_FIFO_blk[16] = 1'b0;
    assign proc_31_data_PIPO_blk[16] = 1'b0;
    assign proc_31_start_FIFO_blk[16] = 1'b0;
    assign proc_31_TLF_FIFO_blk[16] = 1'b0;
    assign proc_31_input_sync_blk[16] = 1'b0;
    assign proc_31_output_sync_blk[16] = 1'b0 | (ap_done_reg_12 & write_back60_U0.ap_done & ~write_back63_U0.ap_done);
    assign proc_dep_vld_vec_31[16] = dl_detect_out ? proc_dep_vld_vec_31_reg[16] : (proc_31_data_FIFO_blk[16] | proc_31_data_PIPO_blk[16] | proc_31_start_FIFO_blk[16] | proc_31_TLF_FIFO_blk[16] | proc_31_input_sync_blk[16] | proc_31_output_sync_blk[16]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_31_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_31_reg <= proc_dep_vld_vec_31;
        end
    end
    assign in_chan_dep_vld_vec_31[0] = dep_chan_vld_0_31;
    assign in_chan_dep_data_vec_31[34 : 0] = dep_chan_data_0_31;
    assign token_in_vec_31[0] = token_0_31;
    assign in_chan_dep_vld_vec_31[1] = dep_chan_vld_15_31;
    assign in_chan_dep_data_vec_31[69 : 35] = dep_chan_data_15_31;
    assign token_in_vec_31[1] = token_15_31;
    assign in_chan_dep_vld_vec_31[2] = dep_chan_vld_19_31;
    assign in_chan_dep_data_vec_31[104 : 70] = dep_chan_data_19_31;
    assign token_in_vec_31[2] = token_19_31;
    assign in_chan_dep_vld_vec_31[3] = dep_chan_vld_20_31;
    assign in_chan_dep_data_vec_31[139 : 105] = dep_chan_data_20_31;
    assign token_in_vec_31[3] = token_20_31;
    assign in_chan_dep_vld_vec_31[4] = dep_chan_vld_21_31;
    assign in_chan_dep_data_vec_31[174 : 140] = dep_chan_data_21_31;
    assign token_in_vec_31[4] = token_21_31;
    assign in_chan_dep_vld_vec_31[5] = dep_chan_vld_22_31;
    assign in_chan_dep_data_vec_31[209 : 175] = dep_chan_data_22_31;
    assign token_in_vec_31[5] = token_22_31;
    assign in_chan_dep_vld_vec_31[6] = dep_chan_vld_23_31;
    assign in_chan_dep_data_vec_31[244 : 210] = dep_chan_data_23_31;
    assign token_in_vec_31[6] = token_23_31;
    assign in_chan_dep_vld_vec_31[7] = dep_chan_vld_24_31;
    assign in_chan_dep_data_vec_31[279 : 245] = dep_chan_data_24_31;
    assign token_in_vec_31[7] = token_24_31;
    assign in_chan_dep_vld_vec_31[8] = dep_chan_vld_25_31;
    assign in_chan_dep_data_vec_31[314 : 280] = dep_chan_data_25_31;
    assign token_in_vec_31[8] = token_25_31;
    assign in_chan_dep_vld_vec_31[9] = dep_chan_vld_26_31;
    assign in_chan_dep_data_vec_31[349 : 315] = dep_chan_data_26_31;
    assign token_in_vec_31[9] = token_26_31;
    assign in_chan_dep_vld_vec_31[10] = dep_chan_vld_27_31;
    assign in_chan_dep_data_vec_31[384 : 350] = dep_chan_data_27_31;
    assign token_in_vec_31[10] = token_27_31;
    assign in_chan_dep_vld_vec_31[11] = dep_chan_vld_28_31;
    assign in_chan_dep_data_vec_31[419 : 385] = dep_chan_data_28_31;
    assign token_in_vec_31[11] = token_28_31;
    assign in_chan_dep_vld_vec_31[12] = dep_chan_vld_29_31;
    assign in_chan_dep_data_vec_31[454 : 420] = dep_chan_data_29_31;
    assign token_in_vec_31[12] = token_29_31;
    assign in_chan_dep_vld_vec_31[13] = dep_chan_vld_30_31;
    assign in_chan_dep_data_vec_31[489 : 455] = dep_chan_data_30_31;
    assign token_in_vec_31[13] = token_30_31;
    assign in_chan_dep_vld_vec_31[14] = dep_chan_vld_32_31;
    assign in_chan_dep_data_vec_31[524 : 490] = dep_chan_data_32_31;
    assign token_in_vec_31[14] = token_32_31;
    assign in_chan_dep_vld_vec_31[15] = dep_chan_vld_33_31;
    assign in_chan_dep_data_vec_31[559 : 525] = dep_chan_data_33_31;
    assign token_in_vec_31[15] = token_33_31;
    assign in_chan_dep_vld_vec_31[16] = dep_chan_vld_34_31;
    assign in_chan_dep_data_vec_31[594 : 560] = dep_chan_data_34_31;
    assign token_in_vec_31[16] = token_34_31;
    assign dep_chan_vld_31_0 = out_chan_dep_vld_vec_31[0];
    assign dep_chan_data_31_0 = out_chan_dep_data_31;
    assign token_31_0 = token_out_vec_31[0];
    assign dep_chan_vld_31_15 = out_chan_dep_vld_vec_31[1];
    assign dep_chan_data_31_15 = out_chan_dep_data_31;
    assign token_31_15 = token_out_vec_31[1];
    assign dep_chan_vld_31_19 = out_chan_dep_vld_vec_31[2];
    assign dep_chan_data_31_19 = out_chan_dep_data_31;
    assign token_31_19 = token_out_vec_31[2];
    assign dep_chan_vld_31_20 = out_chan_dep_vld_vec_31[3];
    assign dep_chan_data_31_20 = out_chan_dep_data_31;
    assign token_31_20 = token_out_vec_31[3];
    assign dep_chan_vld_31_21 = out_chan_dep_vld_vec_31[4];
    assign dep_chan_data_31_21 = out_chan_dep_data_31;
    assign token_31_21 = token_out_vec_31[4];
    assign dep_chan_vld_31_22 = out_chan_dep_vld_vec_31[5];
    assign dep_chan_data_31_22 = out_chan_dep_data_31;
    assign token_31_22 = token_out_vec_31[5];
    assign dep_chan_vld_31_23 = out_chan_dep_vld_vec_31[6];
    assign dep_chan_data_31_23 = out_chan_dep_data_31;
    assign token_31_23 = token_out_vec_31[6];
    assign dep_chan_vld_31_24 = out_chan_dep_vld_vec_31[7];
    assign dep_chan_data_31_24 = out_chan_dep_data_31;
    assign token_31_24 = token_out_vec_31[7];
    assign dep_chan_vld_31_25 = out_chan_dep_vld_vec_31[8];
    assign dep_chan_data_31_25 = out_chan_dep_data_31;
    assign token_31_25 = token_out_vec_31[8];
    assign dep_chan_vld_31_26 = out_chan_dep_vld_vec_31[9];
    assign dep_chan_data_31_26 = out_chan_dep_data_31;
    assign token_31_26 = token_out_vec_31[9];
    assign dep_chan_vld_31_27 = out_chan_dep_vld_vec_31[10];
    assign dep_chan_data_31_27 = out_chan_dep_data_31;
    assign token_31_27 = token_out_vec_31[10];
    assign dep_chan_vld_31_28 = out_chan_dep_vld_vec_31[11];
    assign dep_chan_data_31_28 = out_chan_dep_data_31;
    assign token_31_28 = token_out_vec_31[11];
    assign dep_chan_vld_31_29 = out_chan_dep_vld_vec_31[12];
    assign dep_chan_data_31_29 = out_chan_dep_data_31;
    assign token_31_29 = token_out_vec_31[12];
    assign dep_chan_vld_31_30 = out_chan_dep_vld_vec_31[13];
    assign dep_chan_data_31_30 = out_chan_dep_data_31;
    assign token_31_30 = token_out_vec_31[13];
    assign dep_chan_vld_31_32 = out_chan_dep_vld_vec_31[14];
    assign dep_chan_data_31_32 = out_chan_dep_data_31;
    assign token_31_32 = token_out_vec_31[14];
    assign dep_chan_vld_31_33 = out_chan_dep_vld_vec_31[15];
    assign dep_chan_data_31_33 = out_chan_dep_data_31;
    assign token_31_33 = token_out_vec_31[15];
    assign dep_chan_vld_31_34 = out_chan_dep_vld_vec_31[16];
    assign dep_chan_data_31_34 = out_chan_dep_data_31;
    assign token_31_34 = token_out_vec_31[16];

    // Process: write_back61_U0
    kernel_pr_hls_deadlock_detect_unit #(35, 32, 17, 17) kernel_pr_hls_deadlock_detect_unit_32 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_32),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_32),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_32),
        .token_in_vec(token_in_vec_32),
        .dl_detect_in(dl_detect_out),
        .origin(origin[32]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_32),
        .out_chan_dep_data(out_chan_dep_data_32),
        .token_out_vec(token_out_vec_32),
        .dl_detect_out(dl_in_vec[32]));

    assign proc_32_data_FIFO_blk[0] = 1'b0 | (~write_back61_U0.H_blk_n) | (~write_back61_U0.hyperedge_size_blk_n);
    assign proc_32_data_PIPO_blk[0] = 1'b0;
    assign proc_32_start_FIFO_blk[0] = 1'b0 | (~start_for_write_back61_U0_U.if_empty_n & write_back61_U0.ap_idle & ~start_for_write_back61_U0_U.if_write);
    assign proc_32_TLF_FIFO_blk[0] = 1'b0;
    assign proc_32_input_sync_blk[0] = 1'b0;
    assign proc_32_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_32[0] = dl_detect_out ? proc_dep_vld_vec_32_reg[0] : (proc_32_data_FIFO_blk[0] | proc_32_data_PIPO_blk[0] | proc_32_start_FIFO_blk[0] | proc_32_TLF_FIFO_blk[0] | proc_32_input_sync_blk[0] | proc_32_output_sync_blk[0]);
    assign proc_32_data_FIFO_blk[1] = 1'b0 | (~write_back61_U0.value_stream_V_V13_blk_n);
    assign proc_32_data_PIPO_blk[1] = 1'b0;
    assign proc_32_start_FIFO_blk[1] = 1'b0;
    assign proc_32_TLF_FIFO_blk[1] = 1'b0;
    assign proc_32_input_sync_blk[1] = 1'b0;
    assign proc_32_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_32[1] = dl_detect_out ? proc_dep_vld_vec_32_reg[1] : (proc_32_data_FIFO_blk[1] | proc_32_data_PIPO_blk[1] | proc_32_start_FIFO_blk[1] | proc_32_TLF_FIFO_blk[1] | proc_32_input_sync_blk[1] | proc_32_output_sync_blk[1]);
    assign proc_32_data_FIFO_blk[2] = 1'b0;
    assign proc_32_data_PIPO_blk[2] = 1'b0;
    assign proc_32_start_FIFO_blk[2] = 1'b0;
    assign proc_32_TLF_FIFO_blk[2] = 1'b0;
    assign proc_32_input_sync_blk[2] = 1'b0;
    assign proc_32_output_sync_blk[2] = 1'b0 | (ap_done_reg_13 & write_back61_U0.ap_done & ~write_back48_U0.ap_done);
    assign proc_dep_vld_vec_32[2] = dl_detect_out ? proc_dep_vld_vec_32_reg[2] : (proc_32_data_FIFO_blk[2] | proc_32_data_PIPO_blk[2] | proc_32_start_FIFO_blk[2] | proc_32_TLF_FIFO_blk[2] | proc_32_input_sync_blk[2] | proc_32_output_sync_blk[2]);
    assign proc_32_data_FIFO_blk[3] = 1'b0;
    assign proc_32_data_PIPO_blk[3] = 1'b0;
    assign proc_32_start_FIFO_blk[3] = 1'b0;
    assign proc_32_TLF_FIFO_blk[3] = 1'b0;
    assign proc_32_input_sync_blk[3] = 1'b0;
    assign proc_32_output_sync_blk[3] = 1'b0 | (ap_done_reg_13 & write_back61_U0.ap_done & ~write_back49_U0.ap_done);
    assign proc_dep_vld_vec_32[3] = dl_detect_out ? proc_dep_vld_vec_32_reg[3] : (proc_32_data_FIFO_blk[3] | proc_32_data_PIPO_blk[3] | proc_32_start_FIFO_blk[3] | proc_32_TLF_FIFO_blk[3] | proc_32_input_sync_blk[3] | proc_32_output_sync_blk[3]);
    assign proc_32_data_FIFO_blk[4] = 1'b0;
    assign proc_32_data_PIPO_blk[4] = 1'b0;
    assign proc_32_start_FIFO_blk[4] = 1'b0;
    assign proc_32_TLF_FIFO_blk[4] = 1'b0;
    assign proc_32_input_sync_blk[4] = 1'b0;
    assign proc_32_output_sync_blk[4] = 1'b0 | (ap_done_reg_13 & write_back61_U0.ap_done & ~write_back50_U0.ap_done);
    assign proc_dep_vld_vec_32[4] = dl_detect_out ? proc_dep_vld_vec_32_reg[4] : (proc_32_data_FIFO_blk[4] | proc_32_data_PIPO_blk[4] | proc_32_start_FIFO_blk[4] | proc_32_TLF_FIFO_blk[4] | proc_32_input_sync_blk[4] | proc_32_output_sync_blk[4]);
    assign proc_32_data_FIFO_blk[5] = 1'b0;
    assign proc_32_data_PIPO_blk[5] = 1'b0;
    assign proc_32_start_FIFO_blk[5] = 1'b0;
    assign proc_32_TLF_FIFO_blk[5] = 1'b0;
    assign proc_32_input_sync_blk[5] = 1'b0;
    assign proc_32_output_sync_blk[5] = 1'b0 | (ap_done_reg_13 & write_back61_U0.ap_done & ~write_back51_U0.ap_done);
    assign proc_dep_vld_vec_32[5] = dl_detect_out ? proc_dep_vld_vec_32_reg[5] : (proc_32_data_FIFO_blk[5] | proc_32_data_PIPO_blk[5] | proc_32_start_FIFO_blk[5] | proc_32_TLF_FIFO_blk[5] | proc_32_input_sync_blk[5] | proc_32_output_sync_blk[5]);
    assign proc_32_data_FIFO_blk[6] = 1'b0;
    assign proc_32_data_PIPO_blk[6] = 1'b0;
    assign proc_32_start_FIFO_blk[6] = 1'b0;
    assign proc_32_TLF_FIFO_blk[6] = 1'b0;
    assign proc_32_input_sync_blk[6] = 1'b0;
    assign proc_32_output_sync_blk[6] = 1'b0 | (ap_done_reg_13 & write_back61_U0.ap_done & ~write_back52_U0.ap_done);
    assign proc_dep_vld_vec_32[6] = dl_detect_out ? proc_dep_vld_vec_32_reg[6] : (proc_32_data_FIFO_blk[6] | proc_32_data_PIPO_blk[6] | proc_32_start_FIFO_blk[6] | proc_32_TLF_FIFO_blk[6] | proc_32_input_sync_blk[6] | proc_32_output_sync_blk[6]);
    assign proc_32_data_FIFO_blk[7] = 1'b0;
    assign proc_32_data_PIPO_blk[7] = 1'b0;
    assign proc_32_start_FIFO_blk[7] = 1'b0;
    assign proc_32_TLF_FIFO_blk[7] = 1'b0;
    assign proc_32_input_sync_blk[7] = 1'b0;
    assign proc_32_output_sync_blk[7] = 1'b0 | (ap_done_reg_13 & write_back61_U0.ap_done & ~write_back53_U0.ap_done);
    assign proc_dep_vld_vec_32[7] = dl_detect_out ? proc_dep_vld_vec_32_reg[7] : (proc_32_data_FIFO_blk[7] | proc_32_data_PIPO_blk[7] | proc_32_start_FIFO_blk[7] | proc_32_TLF_FIFO_blk[7] | proc_32_input_sync_blk[7] | proc_32_output_sync_blk[7]);
    assign proc_32_data_FIFO_blk[8] = 1'b0;
    assign proc_32_data_PIPO_blk[8] = 1'b0;
    assign proc_32_start_FIFO_blk[8] = 1'b0;
    assign proc_32_TLF_FIFO_blk[8] = 1'b0;
    assign proc_32_input_sync_blk[8] = 1'b0;
    assign proc_32_output_sync_blk[8] = 1'b0 | (ap_done_reg_13 & write_back61_U0.ap_done & ~write_back54_U0.ap_done);
    assign proc_dep_vld_vec_32[8] = dl_detect_out ? proc_dep_vld_vec_32_reg[8] : (proc_32_data_FIFO_blk[8] | proc_32_data_PIPO_blk[8] | proc_32_start_FIFO_blk[8] | proc_32_TLF_FIFO_blk[8] | proc_32_input_sync_blk[8] | proc_32_output_sync_blk[8]);
    assign proc_32_data_FIFO_blk[9] = 1'b0;
    assign proc_32_data_PIPO_blk[9] = 1'b0;
    assign proc_32_start_FIFO_blk[9] = 1'b0;
    assign proc_32_TLF_FIFO_blk[9] = 1'b0;
    assign proc_32_input_sync_blk[9] = 1'b0;
    assign proc_32_output_sync_blk[9] = 1'b0 | (ap_done_reg_13 & write_back61_U0.ap_done & ~write_back55_U0.ap_done);
    assign proc_dep_vld_vec_32[9] = dl_detect_out ? proc_dep_vld_vec_32_reg[9] : (proc_32_data_FIFO_blk[9] | proc_32_data_PIPO_blk[9] | proc_32_start_FIFO_blk[9] | proc_32_TLF_FIFO_blk[9] | proc_32_input_sync_blk[9] | proc_32_output_sync_blk[9]);
    assign proc_32_data_FIFO_blk[10] = 1'b0;
    assign proc_32_data_PIPO_blk[10] = 1'b0;
    assign proc_32_start_FIFO_blk[10] = 1'b0;
    assign proc_32_TLF_FIFO_blk[10] = 1'b0;
    assign proc_32_input_sync_blk[10] = 1'b0;
    assign proc_32_output_sync_blk[10] = 1'b0 | (ap_done_reg_13 & write_back61_U0.ap_done & ~write_back56_U0.ap_done);
    assign proc_dep_vld_vec_32[10] = dl_detect_out ? proc_dep_vld_vec_32_reg[10] : (proc_32_data_FIFO_blk[10] | proc_32_data_PIPO_blk[10] | proc_32_start_FIFO_blk[10] | proc_32_TLF_FIFO_blk[10] | proc_32_input_sync_blk[10] | proc_32_output_sync_blk[10]);
    assign proc_32_data_FIFO_blk[11] = 1'b0;
    assign proc_32_data_PIPO_blk[11] = 1'b0;
    assign proc_32_start_FIFO_blk[11] = 1'b0;
    assign proc_32_TLF_FIFO_blk[11] = 1'b0;
    assign proc_32_input_sync_blk[11] = 1'b0;
    assign proc_32_output_sync_blk[11] = 1'b0 | (ap_done_reg_13 & write_back61_U0.ap_done & ~write_back57_U0.ap_done);
    assign proc_dep_vld_vec_32[11] = dl_detect_out ? proc_dep_vld_vec_32_reg[11] : (proc_32_data_FIFO_blk[11] | proc_32_data_PIPO_blk[11] | proc_32_start_FIFO_blk[11] | proc_32_TLF_FIFO_blk[11] | proc_32_input_sync_blk[11] | proc_32_output_sync_blk[11]);
    assign proc_32_data_FIFO_blk[12] = 1'b0;
    assign proc_32_data_PIPO_blk[12] = 1'b0;
    assign proc_32_start_FIFO_blk[12] = 1'b0;
    assign proc_32_TLF_FIFO_blk[12] = 1'b0;
    assign proc_32_input_sync_blk[12] = 1'b0;
    assign proc_32_output_sync_blk[12] = 1'b0 | (ap_done_reg_13 & write_back61_U0.ap_done & ~write_back58_U0.ap_done);
    assign proc_dep_vld_vec_32[12] = dl_detect_out ? proc_dep_vld_vec_32_reg[12] : (proc_32_data_FIFO_blk[12] | proc_32_data_PIPO_blk[12] | proc_32_start_FIFO_blk[12] | proc_32_TLF_FIFO_blk[12] | proc_32_input_sync_blk[12] | proc_32_output_sync_blk[12]);
    assign proc_32_data_FIFO_blk[13] = 1'b0;
    assign proc_32_data_PIPO_blk[13] = 1'b0;
    assign proc_32_start_FIFO_blk[13] = 1'b0;
    assign proc_32_TLF_FIFO_blk[13] = 1'b0;
    assign proc_32_input_sync_blk[13] = 1'b0;
    assign proc_32_output_sync_blk[13] = 1'b0 | (ap_done_reg_13 & write_back61_U0.ap_done & ~write_back59_U0.ap_done);
    assign proc_dep_vld_vec_32[13] = dl_detect_out ? proc_dep_vld_vec_32_reg[13] : (proc_32_data_FIFO_blk[13] | proc_32_data_PIPO_blk[13] | proc_32_start_FIFO_blk[13] | proc_32_TLF_FIFO_blk[13] | proc_32_input_sync_blk[13] | proc_32_output_sync_blk[13]);
    assign proc_32_data_FIFO_blk[14] = 1'b0;
    assign proc_32_data_PIPO_blk[14] = 1'b0;
    assign proc_32_start_FIFO_blk[14] = 1'b0;
    assign proc_32_TLF_FIFO_blk[14] = 1'b0;
    assign proc_32_input_sync_blk[14] = 1'b0;
    assign proc_32_output_sync_blk[14] = 1'b0 | (ap_done_reg_13 & write_back61_U0.ap_done & ~write_back60_U0.ap_done);
    assign proc_dep_vld_vec_32[14] = dl_detect_out ? proc_dep_vld_vec_32_reg[14] : (proc_32_data_FIFO_blk[14] | proc_32_data_PIPO_blk[14] | proc_32_start_FIFO_blk[14] | proc_32_TLF_FIFO_blk[14] | proc_32_input_sync_blk[14] | proc_32_output_sync_blk[14]);
    assign proc_32_data_FIFO_blk[15] = 1'b0;
    assign proc_32_data_PIPO_blk[15] = 1'b0;
    assign proc_32_start_FIFO_blk[15] = 1'b0;
    assign proc_32_TLF_FIFO_blk[15] = 1'b0;
    assign proc_32_input_sync_blk[15] = 1'b0;
    assign proc_32_output_sync_blk[15] = 1'b0 | (ap_done_reg_13 & write_back61_U0.ap_done & ~write_back62_U0.ap_done);
    assign proc_dep_vld_vec_32[15] = dl_detect_out ? proc_dep_vld_vec_32_reg[15] : (proc_32_data_FIFO_blk[15] | proc_32_data_PIPO_blk[15] | proc_32_start_FIFO_blk[15] | proc_32_TLF_FIFO_blk[15] | proc_32_input_sync_blk[15] | proc_32_output_sync_blk[15]);
    assign proc_32_data_FIFO_blk[16] = 1'b0;
    assign proc_32_data_PIPO_blk[16] = 1'b0;
    assign proc_32_start_FIFO_blk[16] = 1'b0;
    assign proc_32_TLF_FIFO_blk[16] = 1'b0;
    assign proc_32_input_sync_blk[16] = 1'b0;
    assign proc_32_output_sync_blk[16] = 1'b0 | (ap_done_reg_13 & write_back61_U0.ap_done & ~write_back63_U0.ap_done);
    assign proc_dep_vld_vec_32[16] = dl_detect_out ? proc_dep_vld_vec_32_reg[16] : (proc_32_data_FIFO_blk[16] | proc_32_data_PIPO_blk[16] | proc_32_start_FIFO_blk[16] | proc_32_TLF_FIFO_blk[16] | proc_32_input_sync_blk[16] | proc_32_output_sync_blk[16]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_32_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_32_reg <= proc_dep_vld_vec_32;
        end
    end
    assign in_chan_dep_vld_vec_32[0] = dep_chan_vld_0_32;
    assign in_chan_dep_data_vec_32[34 : 0] = dep_chan_data_0_32;
    assign token_in_vec_32[0] = token_0_32;
    assign in_chan_dep_vld_vec_32[1] = dep_chan_vld_16_32;
    assign in_chan_dep_data_vec_32[69 : 35] = dep_chan_data_16_32;
    assign token_in_vec_32[1] = token_16_32;
    assign in_chan_dep_vld_vec_32[2] = dep_chan_vld_19_32;
    assign in_chan_dep_data_vec_32[104 : 70] = dep_chan_data_19_32;
    assign token_in_vec_32[2] = token_19_32;
    assign in_chan_dep_vld_vec_32[3] = dep_chan_vld_20_32;
    assign in_chan_dep_data_vec_32[139 : 105] = dep_chan_data_20_32;
    assign token_in_vec_32[3] = token_20_32;
    assign in_chan_dep_vld_vec_32[4] = dep_chan_vld_21_32;
    assign in_chan_dep_data_vec_32[174 : 140] = dep_chan_data_21_32;
    assign token_in_vec_32[4] = token_21_32;
    assign in_chan_dep_vld_vec_32[5] = dep_chan_vld_22_32;
    assign in_chan_dep_data_vec_32[209 : 175] = dep_chan_data_22_32;
    assign token_in_vec_32[5] = token_22_32;
    assign in_chan_dep_vld_vec_32[6] = dep_chan_vld_23_32;
    assign in_chan_dep_data_vec_32[244 : 210] = dep_chan_data_23_32;
    assign token_in_vec_32[6] = token_23_32;
    assign in_chan_dep_vld_vec_32[7] = dep_chan_vld_24_32;
    assign in_chan_dep_data_vec_32[279 : 245] = dep_chan_data_24_32;
    assign token_in_vec_32[7] = token_24_32;
    assign in_chan_dep_vld_vec_32[8] = dep_chan_vld_25_32;
    assign in_chan_dep_data_vec_32[314 : 280] = dep_chan_data_25_32;
    assign token_in_vec_32[8] = token_25_32;
    assign in_chan_dep_vld_vec_32[9] = dep_chan_vld_26_32;
    assign in_chan_dep_data_vec_32[349 : 315] = dep_chan_data_26_32;
    assign token_in_vec_32[9] = token_26_32;
    assign in_chan_dep_vld_vec_32[10] = dep_chan_vld_27_32;
    assign in_chan_dep_data_vec_32[384 : 350] = dep_chan_data_27_32;
    assign token_in_vec_32[10] = token_27_32;
    assign in_chan_dep_vld_vec_32[11] = dep_chan_vld_28_32;
    assign in_chan_dep_data_vec_32[419 : 385] = dep_chan_data_28_32;
    assign token_in_vec_32[11] = token_28_32;
    assign in_chan_dep_vld_vec_32[12] = dep_chan_vld_29_32;
    assign in_chan_dep_data_vec_32[454 : 420] = dep_chan_data_29_32;
    assign token_in_vec_32[12] = token_29_32;
    assign in_chan_dep_vld_vec_32[13] = dep_chan_vld_30_32;
    assign in_chan_dep_data_vec_32[489 : 455] = dep_chan_data_30_32;
    assign token_in_vec_32[13] = token_30_32;
    assign in_chan_dep_vld_vec_32[14] = dep_chan_vld_31_32;
    assign in_chan_dep_data_vec_32[524 : 490] = dep_chan_data_31_32;
    assign token_in_vec_32[14] = token_31_32;
    assign in_chan_dep_vld_vec_32[15] = dep_chan_vld_33_32;
    assign in_chan_dep_data_vec_32[559 : 525] = dep_chan_data_33_32;
    assign token_in_vec_32[15] = token_33_32;
    assign in_chan_dep_vld_vec_32[16] = dep_chan_vld_34_32;
    assign in_chan_dep_data_vec_32[594 : 560] = dep_chan_data_34_32;
    assign token_in_vec_32[16] = token_34_32;
    assign dep_chan_vld_32_0 = out_chan_dep_vld_vec_32[0];
    assign dep_chan_data_32_0 = out_chan_dep_data_32;
    assign token_32_0 = token_out_vec_32[0];
    assign dep_chan_vld_32_16 = out_chan_dep_vld_vec_32[1];
    assign dep_chan_data_32_16 = out_chan_dep_data_32;
    assign token_32_16 = token_out_vec_32[1];
    assign dep_chan_vld_32_19 = out_chan_dep_vld_vec_32[2];
    assign dep_chan_data_32_19 = out_chan_dep_data_32;
    assign token_32_19 = token_out_vec_32[2];
    assign dep_chan_vld_32_20 = out_chan_dep_vld_vec_32[3];
    assign dep_chan_data_32_20 = out_chan_dep_data_32;
    assign token_32_20 = token_out_vec_32[3];
    assign dep_chan_vld_32_21 = out_chan_dep_vld_vec_32[4];
    assign dep_chan_data_32_21 = out_chan_dep_data_32;
    assign token_32_21 = token_out_vec_32[4];
    assign dep_chan_vld_32_22 = out_chan_dep_vld_vec_32[5];
    assign dep_chan_data_32_22 = out_chan_dep_data_32;
    assign token_32_22 = token_out_vec_32[5];
    assign dep_chan_vld_32_23 = out_chan_dep_vld_vec_32[6];
    assign dep_chan_data_32_23 = out_chan_dep_data_32;
    assign token_32_23 = token_out_vec_32[6];
    assign dep_chan_vld_32_24 = out_chan_dep_vld_vec_32[7];
    assign dep_chan_data_32_24 = out_chan_dep_data_32;
    assign token_32_24 = token_out_vec_32[7];
    assign dep_chan_vld_32_25 = out_chan_dep_vld_vec_32[8];
    assign dep_chan_data_32_25 = out_chan_dep_data_32;
    assign token_32_25 = token_out_vec_32[8];
    assign dep_chan_vld_32_26 = out_chan_dep_vld_vec_32[9];
    assign dep_chan_data_32_26 = out_chan_dep_data_32;
    assign token_32_26 = token_out_vec_32[9];
    assign dep_chan_vld_32_27 = out_chan_dep_vld_vec_32[10];
    assign dep_chan_data_32_27 = out_chan_dep_data_32;
    assign token_32_27 = token_out_vec_32[10];
    assign dep_chan_vld_32_28 = out_chan_dep_vld_vec_32[11];
    assign dep_chan_data_32_28 = out_chan_dep_data_32;
    assign token_32_28 = token_out_vec_32[11];
    assign dep_chan_vld_32_29 = out_chan_dep_vld_vec_32[12];
    assign dep_chan_data_32_29 = out_chan_dep_data_32;
    assign token_32_29 = token_out_vec_32[12];
    assign dep_chan_vld_32_30 = out_chan_dep_vld_vec_32[13];
    assign dep_chan_data_32_30 = out_chan_dep_data_32;
    assign token_32_30 = token_out_vec_32[13];
    assign dep_chan_vld_32_31 = out_chan_dep_vld_vec_32[14];
    assign dep_chan_data_32_31 = out_chan_dep_data_32;
    assign token_32_31 = token_out_vec_32[14];
    assign dep_chan_vld_32_33 = out_chan_dep_vld_vec_32[15];
    assign dep_chan_data_32_33 = out_chan_dep_data_32;
    assign token_32_33 = token_out_vec_32[15];
    assign dep_chan_vld_32_34 = out_chan_dep_vld_vec_32[16];
    assign dep_chan_data_32_34 = out_chan_dep_data_32;
    assign token_32_34 = token_out_vec_32[16];

    // Process: write_back62_U0
    kernel_pr_hls_deadlock_detect_unit #(35, 33, 17, 17) kernel_pr_hls_deadlock_detect_unit_33 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_33),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_33),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_33),
        .token_in_vec(token_in_vec_33),
        .dl_detect_in(dl_detect_out),
        .origin(origin[33]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_33),
        .out_chan_dep_data(out_chan_dep_data_33),
        .token_out_vec(token_out_vec_33),
        .dl_detect_out(dl_in_vec[33]));

    assign proc_33_data_FIFO_blk[0] = 1'b0 | (~write_back62_U0.H_blk_n) | (~write_back62_U0.hyperedge_size_blk_n);
    assign proc_33_data_PIPO_blk[0] = 1'b0;
    assign proc_33_start_FIFO_blk[0] = 1'b0 | (~start_for_write_back62_U0_U.if_empty_n & write_back62_U0.ap_idle & ~start_for_write_back62_U0_U.if_write);
    assign proc_33_TLF_FIFO_blk[0] = 1'b0;
    assign proc_33_input_sync_blk[0] = 1'b0;
    assign proc_33_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_33[0] = dl_detect_out ? proc_dep_vld_vec_33_reg[0] : (proc_33_data_FIFO_blk[0] | proc_33_data_PIPO_blk[0] | proc_33_start_FIFO_blk[0] | proc_33_TLF_FIFO_blk[0] | proc_33_input_sync_blk[0] | proc_33_output_sync_blk[0]);
    assign proc_33_data_FIFO_blk[1] = 1'b0 | (~write_back62_U0.value_stream_V_V14_blk_n);
    assign proc_33_data_PIPO_blk[1] = 1'b0;
    assign proc_33_start_FIFO_blk[1] = 1'b0;
    assign proc_33_TLF_FIFO_blk[1] = 1'b0;
    assign proc_33_input_sync_blk[1] = 1'b0;
    assign proc_33_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_33[1] = dl_detect_out ? proc_dep_vld_vec_33_reg[1] : (proc_33_data_FIFO_blk[1] | proc_33_data_PIPO_blk[1] | proc_33_start_FIFO_blk[1] | proc_33_TLF_FIFO_blk[1] | proc_33_input_sync_blk[1] | proc_33_output_sync_blk[1]);
    assign proc_33_data_FIFO_blk[2] = 1'b0;
    assign proc_33_data_PIPO_blk[2] = 1'b0;
    assign proc_33_start_FIFO_blk[2] = 1'b0;
    assign proc_33_TLF_FIFO_blk[2] = 1'b0;
    assign proc_33_input_sync_blk[2] = 1'b0;
    assign proc_33_output_sync_blk[2] = 1'b0 | (ap_done_reg_14 & write_back62_U0.ap_done & ~write_back48_U0.ap_done);
    assign proc_dep_vld_vec_33[2] = dl_detect_out ? proc_dep_vld_vec_33_reg[2] : (proc_33_data_FIFO_blk[2] | proc_33_data_PIPO_blk[2] | proc_33_start_FIFO_blk[2] | proc_33_TLF_FIFO_blk[2] | proc_33_input_sync_blk[2] | proc_33_output_sync_blk[2]);
    assign proc_33_data_FIFO_blk[3] = 1'b0;
    assign proc_33_data_PIPO_blk[3] = 1'b0;
    assign proc_33_start_FIFO_blk[3] = 1'b0;
    assign proc_33_TLF_FIFO_blk[3] = 1'b0;
    assign proc_33_input_sync_blk[3] = 1'b0;
    assign proc_33_output_sync_blk[3] = 1'b0 | (ap_done_reg_14 & write_back62_U0.ap_done & ~write_back49_U0.ap_done);
    assign proc_dep_vld_vec_33[3] = dl_detect_out ? proc_dep_vld_vec_33_reg[3] : (proc_33_data_FIFO_blk[3] | proc_33_data_PIPO_blk[3] | proc_33_start_FIFO_blk[3] | proc_33_TLF_FIFO_blk[3] | proc_33_input_sync_blk[3] | proc_33_output_sync_blk[3]);
    assign proc_33_data_FIFO_blk[4] = 1'b0;
    assign proc_33_data_PIPO_blk[4] = 1'b0;
    assign proc_33_start_FIFO_blk[4] = 1'b0;
    assign proc_33_TLF_FIFO_blk[4] = 1'b0;
    assign proc_33_input_sync_blk[4] = 1'b0;
    assign proc_33_output_sync_blk[4] = 1'b0 | (ap_done_reg_14 & write_back62_U0.ap_done & ~write_back50_U0.ap_done);
    assign proc_dep_vld_vec_33[4] = dl_detect_out ? proc_dep_vld_vec_33_reg[4] : (proc_33_data_FIFO_blk[4] | proc_33_data_PIPO_blk[4] | proc_33_start_FIFO_blk[4] | proc_33_TLF_FIFO_blk[4] | proc_33_input_sync_blk[4] | proc_33_output_sync_blk[4]);
    assign proc_33_data_FIFO_blk[5] = 1'b0;
    assign proc_33_data_PIPO_blk[5] = 1'b0;
    assign proc_33_start_FIFO_blk[5] = 1'b0;
    assign proc_33_TLF_FIFO_blk[5] = 1'b0;
    assign proc_33_input_sync_blk[5] = 1'b0;
    assign proc_33_output_sync_blk[5] = 1'b0 | (ap_done_reg_14 & write_back62_U0.ap_done & ~write_back51_U0.ap_done);
    assign proc_dep_vld_vec_33[5] = dl_detect_out ? proc_dep_vld_vec_33_reg[5] : (proc_33_data_FIFO_blk[5] | proc_33_data_PIPO_blk[5] | proc_33_start_FIFO_blk[5] | proc_33_TLF_FIFO_blk[5] | proc_33_input_sync_blk[5] | proc_33_output_sync_blk[5]);
    assign proc_33_data_FIFO_blk[6] = 1'b0;
    assign proc_33_data_PIPO_blk[6] = 1'b0;
    assign proc_33_start_FIFO_blk[6] = 1'b0;
    assign proc_33_TLF_FIFO_blk[6] = 1'b0;
    assign proc_33_input_sync_blk[6] = 1'b0;
    assign proc_33_output_sync_blk[6] = 1'b0 | (ap_done_reg_14 & write_back62_U0.ap_done & ~write_back52_U0.ap_done);
    assign proc_dep_vld_vec_33[6] = dl_detect_out ? proc_dep_vld_vec_33_reg[6] : (proc_33_data_FIFO_blk[6] | proc_33_data_PIPO_blk[6] | proc_33_start_FIFO_blk[6] | proc_33_TLF_FIFO_blk[6] | proc_33_input_sync_blk[6] | proc_33_output_sync_blk[6]);
    assign proc_33_data_FIFO_blk[7] = 1'b0;
    assign proc_33_data_PIPO_blk[7] = 1'b0;
    assign proc_33_start_FIFO_blk[7] = 1'b0;
    assign proc_33_TLF_FIFO_blk[7] = 1'b0;
    assign proc_33_input_sync_blk[7] = 1'b0;
    assign proc_33_output_sync_blk[7] = 1'b0 | (ap_done_reg_14 & write_back62_U0.ap_done & ~write_back53_U0.ap_done);
    assign proc_dep_vld_vec_33[7] = dl_detect_out ? proc_dep_vld_vec_33_reg[7] : (proc_33_data_FIFO_blk[7] | proc_33_data_PIPO_blk[7] | proc_33_start_FIFO_blk[7] | proc_33_TLF_FIFO_blk[7] | proc_33_input_sync_blk[7] | proc_33_output_sync_blk[7]);
    assign proc_33_data_FIFO_blk[8] = 1'b0;
    assign proc_33_data_PIPO_blk[8] = 1'b0;
    assign proc_33_start_FIFO_blk[8] = 1'b0;
    assign proc_33_TLF_FIFO_blk[8] = 1'b0;
    assign proc_33_input_sync_blk[8] = 1'b0;
    assign proc_33_output_sync_blk[8] = 1'b0 | (ap_done_reg_14 & write_back62_U0.ap_done & ~write_back54_U0.ap_done);
    assign proc_dep_vld_vec_33[8] = dl_detect_out ? proc_dep_vld_vec_33_reg[8] : (proc_33_data_FIFO_blk[8] | proc_33_data_PIPO_blk[8] | proc_33_start_FIFO_blk[8] | proc_33_TLF_FIFO_blk[8] | proc_33_input_sync_blk[8] | proc_33_output_sync_blk[8]);
    assign proc_33_data_FIFO_blk[9] = 1'b0;
    assign proc_33_data_PIPO_blk[9] = 1'b0;
    assign proc_33_start_FIFO_blk[9] = 1'b0;
    assign proc_33_TLF_FIFO_blk[9] = 1'b0;
    assign proc_33_input_sync_blk[9] = 1'b0;
    assign proc_33_output_sync_blk[9] = 1'b0 | (ap_done_reg_14 & write_back62_U0.ap_done & ~write_back55_U0.ap_done);
    assign proc_dep_vld_vec_33[9] = dl_detect_out ? proc_dep_vld_vec_33_reg[9] : (proc_33_data_FIFO_blk[9] | proc_33_data_PIPO_blk[9] | proc_33_start_FIFO_blk[9] | proc_33_TLF_FIFO_blk[9] | proc_33_input_sync_blk[9] | proc_33_output_sync_blk[9]);
    assign proc_33_data_FIFO_blk[10] = 1'b0;
    assign proc_33_data_PIPO_blk[10] = 1'b0;
    assign proc_33_start_FIFO_blk[10] = 1'b0;
    assign proc_33_TLF_FIFO_blk[10] = 1'b0;
    assign proc_33_input_sync_blk[10] = 1'b0;
    assign proc_33_output_sync_blk[10] = 1'b0 | (ap_done_reg_14 & write_back62_U0.ap_done & ~write_back56_U0.ap_done);
    assign proc_dep_vld_vec_33[10] = dl_detect_out ? proc_dep_vld_vec_33_reg[10] : (proc_33_data_FIFO_blk[10] | proc_33_data_PIPO_blk[10] | proc_33_start_FIFO_blk[10] | proc_33_TLF_FIFO_blk[10] | proc_33_input_sync_blk[10] | proc_33_output_sync_blk[10]);
    assign proc_33_data_FIFO_blk[11] = 1'b0;
    assign proc_33_data_PIPO_blk[11] = 1'b0;
    assign proc_33_start_FIFO_blk[11] = 1'b0;
    assign proc_33_TLF_FIFO_blk[11] = 1'b0;
    assign proc_33_input_sync_blk[11] = 1'b0;
    assign proc_33_output_sync_blk[11] = 1'b0 | (ap_done_reg_14 & write_back62_U0.ap_done & ~write_back57_U0.ap_done);
    assign proc_dep_vld_vec_33[11] = dl_detect_out ? proc_dep_vld_vec_33_reg[11] : (proc_33_data_FIFO_blk[11] | proc_33_data_PIPO_blk[11] | proc_33_start_FIFO_blk[11] | proc_33_TLF_FIFO_blk[11] | proc_33_input_sync_blk[11] | proc_33_output_sync_blk[11]);
    assign proc_33_data_FIFO_blk[12] = 1'b0;
    assign proc_33_data_PIPO_blk[12] = 1'b0;
    assign proc_33_start_FIFO_blk[12] = 1'b0;
    assign proc_33_TLF_FIFO_blk[12] = 1'b0;
    assign proc_33_input_sync_blk[12] = 1'b0;
    assign proc_33_output_sync_blk[12] = 1'b0 | (ap_done_reg_14 & write_back62_U0.ap_done & ~write_back58_U0.ap_done);
    assign proc_dep_vld_vec_33[12] = dl_detect_out ? proc_dep_vld_vec_33_reg[12] : (proc_33_data_FIFO_blk[12] | proc_33_data_PIPO_blk[12] | proc_33_start_FIFO_blk[12] | proc_33_TLF_FIFO_blk[12] | proc_33_input_sync_blk[12] | proc_33_output_sync_blk[12]);
    assign proc_33_data_FIFO_blk[13] = 1'b0;
    assign proc_33_data_PIPO_blk[13] = 1'b0;
    assign proc_33_start_FIFO_blk[13] = 1'b0;
    assign proc_33_TLF_FIFO_blk[13] = 1'b0;
    assign proc_33_input_sync_blk[13] = 1'b0;
    assign proc_33_output_sync_blk[13] = 1'b0 | (ap_done_reg_14 & write_back62_U0.ap_done & ~write_back59_U0.ap_done);
    assign proc_dep_vld_vec_33[13] = dl_detect_out ? proc_dep_vld_vec_33_reg[13] : (proc_33_data_FIFO_blk[13] | proc_33_data_PIPO_blk[13] | proc_33_start_FIFO_blk[13] | proc_33_TLF_FIFO_blk[13] | proc_33_input_sync_blk[13] | proc_33_output_sync_blk[13]);
    assign proc_33_data_FIFO_blk[14] = 1'b0;
    assign proc_33_data_PIPO_blk[14] = 1'b0;
    assign proc_33_start_FIFO_blk[14] = 1'b0;
    assign proc_33_TLF_FIFO_blk[14] = 1'b0;
    assign proc_33_input_sync_blk[14] = 1'b0;
    assign proc_33_output_sync_blk[14] = 1'b0 | (ap_done_reg_14 & write_back62_U0.ap_done & ~write_back60_U0.ap_done);
    assign proc_dep_vld_vec_33[14] = dl_detect_out ? proc_dep_vld_vec_33_reg[14] : (proc_33_data_FIFO_blk[14] | proc_33_data_PIPO_blk[14] | proc_33_start_FIFO_blk[14] | proc_33_TLF_FIFO_blk[14] | proc_33_input_sync_blk[14] | proc_33_output_sync_blk[14]);
    assign proc_33_data_FIFO_blk[15] = 1'b0;
    assign proc_33_data_PIPO_blk[15] = 1'b0;
    assign proc_33_start_FIFO_blk[15] = 1'b0;
    assign proc_33_TLF_FIFO_blk[15] = 1'b0;
    assign proc_33_input_sync_blk[15] = 1'b0;
    assign proc_33_output_sync_blk[15] = 1'b0 | (ap_done_reg_14 & write_back62_U0.ap_done & ~write_back61_U0.ap_done);
    assign proc_dep_vld_vec_33[15] = dl_detect_out ? proc_dep_vld_vec_33_reg[15] : (proc_33_data_FIFO_blk[15] | proc_33_data_PIPO_blk[15] | proc_33_start_FIFO_blk[15] | proc_33_TLF_FIFO_blk[15] | proc_33_input_sync_blk[15] | proc_33_output_sync_blk[15]);
    assign proc_33_data_FIFO_blk[16] = 1'b0;
    assign proc_33_data_PIPO_blk[16] = 1'b0;
    assign proc_33_start_FIFO_blk[16] = 1'b0;
    assign proc_33_TLF_FIFO_blk[16] = 1'b0;
    assign proc_33_input_sync_blk[16] = 1'b0;
    assign proc_33_output_sync_blk[16] = 1'b0 | (ap_done_reg_14 & write_back62_U0.ap_done & ~write_back63_U0.ap_done);
    assign proc_dep_vld_vec_33[16] = dl_detect_out ? proc_dep_vld_vec_33_reg[16] : (proc_33_data_FIFO_blk[16] | proc_33_data_PIPO_blk[16] | proc_33_start_FIFO_blk[16] | proc_33_TLF_FIFO_blk[16] | proc_33_input_sync_blk[16] | proc_33_output_sync_blk[16]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_33_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_33_reg <= proc_dep_vld_vec_33;
        end
    end
    assign in_chan_dep_vld_vec_33[0] = dep_chan_vld_0_33;
    assign in_chan_dep_data_vec_33[34 : 0] = dep_chan_data_0_33;
    assign token_in_vec_33[0] = token_0_33;
    assign in_chan_dep_vld_vec_33[1] = dep_chan_vld_17_33;
    assign in_chan_dep_data_vec_33[69 : 35] = dep_chan_data_17_33;
    assign token_in_vec_33[1] = token_17_33;
    assign in_chan_dep_vld_vec_33[2] = dep_chan_vld_19_33;
    assign in_chan_dep_data_vec_33[104 : 70] = dep_chan_data_19_33;
    assign token_in_vec_33[2] = token_19_33;
    assign in_chan_dep_vld_vec_33[3] = dep_chan_vld_20_33;
    assign in_chan_dep_data_vec_33[139 : 105] = dep_chan_data_20_33;
    assign token_in_vec_33[3] = token_20_33;
    assign in_chan_dep_vld_vec_33[4] = dep_chan_vld_21_33;
    assign in_chan_dep_data_vec_33[174 : 140] = dep_chan_data_21_33;
    assign token_in_vec_33[4] = token_21_33;
    assign in_chan_dep_vld_vec_33[5] = dep_chan_vld_22_33;
    assign in_chan_dep_data_vec_33[209 : 175] = dep_chan_data_22_33;
    assign token_in_vec_33[5] = token_22_33;
    assign in_chan_dep_vld_vec_33[6] = dep_chan_vld_23_33;
    assign in_chan_dep_data_vec_33[244 : 210] = dep_chan_data_23_33;
    assign token_in_vec_33[6] = token_23_33;
    assign in_chan_dep_vld_vec_33[7] = dep_chan_vld_24_33;
    assign in_chan_dep_data_vec_33[279 : 245] = dep_chan_data_24_33;
    assign token_in_vec_33[7] = token_24_33;
    assign in_chan_dep_vld_vec_33[8] = dep_chan_vld_25_33;
    assign in_chan_dep_data_vec_33[314 : 280] = dep_chan_data_25_33;
    assign token_in_vec_33[8] = token_25_33;
    assign in_chan_dep_vld_vec_33[9] = dep_chan_vld_26_33;
    assign in_chan_dep_data_vec_33[349 : 315] = dep_chan_data_26_33;
    assign token_in_vec_33[9] = token_26_33;
    assign in_chan_dep_vld_vec_33[10] = dep_chan_vld_27_33;
    assign in_chan_dep_data_vec_33[384 : 350] = dep_chan_data_27_33;
    assign token_in_vec_33[10] = token_27_33;
    assign in_chan_dep_vld_vec_33[11] = dep_chan_vld_28_33;
    assign in_chan_dep_data_vec_33[419 : 385] = dep_chan_data_28_33;
    assign token_in_vec_33[11] = token_28_33;
    assign in_chan_dep_vld_vec_33[12] = dep_chan_vld_29_33;
    assign in_chan_dep_data_vec_33[454 : 420] = dep_chan_data_29_33;
    assign token_in_vec_33[12] = token_29_33;
    assign in_chan_dep_vld_vec_33[13] = dep_chan_vld_30_33;
    assign in_chan_dep_data_vec_33[489 : 455] = dep_chan_data_30_33;
    assign token_in_vec_33[13] = token_30_33;
    assign in_chan_dep_vld_vec_33[14] = dep_chan_vld_31_33;
    assign in_chan_dep_data_vec_33[524 : 490] = dep_chan_data_31_33;
    assign token_in_vec_33[14] = token_31_33;
    assign in_chan_dep_vld_vec_33[15] = dep_chan_vld_32_33;
    assign in_chan_dep_data_vec_33[559 : 525] = dep_chan_data_32_33;
    assign token_in_vec_33[15] = token_32_33;
    assign in_chan_dep_vld_vec_33[16] = dep_chan_vld_34_33;
    assign in_chan_dep_data_vec_33[594 : 560] = dep_chan_data_34_33;
    assign token_in_vec_33[16] = token_34_33;
    assign dep_chan_vld_33_0 = out_chan_dep_vld_vec_33[0];
    assign dep_chan_data_33_0 = out_chan_dep_data_33;
    assign token_33_0 = token_out_vec_33[0];
    assign dep_chan_vld_33_17 = out_chan_dep_vld_vec_33[1];
    assign dep_chan_data_33_17 = out_chan_dep_data_33;
    assign token_33_17 = token_out_vec_33[1];
    assign dep_chan_vld_33_19 = out_chan_dep_vld_vec_33[2];
    assign dep_chan_data_33_19 = out_chan_dep_data_33;
    assign token_33_19 = token_out_vec_33[2];
    assign dep_chan_vld_33_20 = out_chan_dep_vld_vec_33[3];
    assign dep_chan_data_33_20 = out_chan_dep_data_33;
    assign token_33_20 = token_out_vec_33[3];
    assign dep_chan_vld_33_21 = out_chan_dep_vld_vec_33[4];
    assign dep_chan_data_33_21 = out_chan_dep_data_33;
    assign token_33_21 = token_out_vec_33[4];
    assign dep_chan_vld_33_22 = out_chan_dep_vld_vec_33[5];
    assign dep_chan_data_33_22 = out_chan_dep_data_33;
    assign token_33_22 = token_out_vec_33[5];
    assign dep_chan_vld_33_23 = out_chan_dep_vld_vec_33[6];
    assign dep_chan_data_33_23 = out_chan_dep_data_33;
    assign token_33_23 = token_out_vec_33[6];
    assign dep_chan_vld_33_24 = out_chan_dep_vld_vec_33[7];
    assign dep_chan_data_33_24 = out_chan_dep_data_33;
    assign token_33_24 = token_out_vec_33[7];
    assign dep_chan_vld_33_25 = out_chan_dep_vld_vec_33[8];
    assign dep_chan_data_33_25 = out_chan_dep_data_33;
    assign token_33_25 = token_out_vec_33[8];
    assign dep_chan_vld_33_26 = out_chan_dep_vld_vec_33[9];
    assign dep_chan_data_33_26 = out_chan_dep_data_33;
    assign token_33_26 = token_out_vec_33[9];
    assign dep_chan_vld_33_27 = out_chan_dep_vld_vec_33[10];
    assign dep_chan_data_33_27 = out_chan_dep_data_33;
    assign token_33_27 = token_out_vec_33[10];
    assign dep_chan_vld_33_28 = out_chan_dep_vld_vec_33[11];
    assign dep_chan_data_33_28 = out_chan_dep_data_33;
    assign token_33_28 = token_out_vec_33[11];
    assign dep_chan_vld_33_29 = out_chan_dep_vld_vec_33[12];
    assign dep_chan_data_33_29 = out_chan_dep_data_33;
    assign token_33_29 = token_out_vec_33[12];
    assign dep_chan_vld_33_30 = out_chan_dep_vld_vec_33[13];
    assign dep_chan_data_33_30 = out_chan_dep_data_33;
    assign token_33_30 = token_out_vec_33[13];
    assign dep_chan_vld_33_31 = out_chan_dep_vld_vec_33[14];
    assign dep_chan_data_33_31 = out_chan_dep_data_33;
    assign token_33_31 = token_out_vec_33[14];
    assign dep_chan_vld_33_32 = out_chan_dep_vld_vec_33[15];
    assign dep_chan_data_33_32 = out_chan_dep_data_33;
    assign token_33_32 = token_out_vec_33[15];
    assign dep_chan_vld_33_34 = out_chan_dep_vld_vec_33[16];
    assign dep_chan_data_33_34 = out_chan_dep_data_33;
    assign token_33_34 = token_out_vec_33[16];

    // Process: write_back63_U0
    kernel_pr_hls_deadlock_detect_unit #(35, 34, 17, 17) kernel_pr_hls_deadlock_detect_unit_34 (
        .reset(reset),
        .clock(clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_34),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_34),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_34),
        .token_in_vec(token_in_vec_34),
        .dl_detect_in(dl_detect_out),
        .origin(origin[34]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_34),
        .out_chan_dep_data(out_chan_dep_data_34),
        .token_out_vec(token_out_vec_34),
        .dl_detect_out(dl_in_vec[34]));

    assign proc_34_data_FIFO_blk[0] = 1'b0 | (~write_back63_U0.H_blk_n) | (~write_back63_U0.hyperedge_size_blk_n);
    assign proc_34_data_PIPO_blk[0] = 1'b0;
    assign proc_34_start_FIFO_blk[0] = 1'b0 | (~start_for_write_back63_U0_U.if_empty_n & write_back63_U0.ap_idle & ~start_for_write_back63_U0_U.if_write);
    assign proc_34_TLF_FIFO_blk[0] = 1'b0;
    assign proc_34_input_sync_blk[0] = 1'b0;
    assign proc_34_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_34[0] = dl_detect_out ? proc_dep_vld_vec_34_reg[0] : (proc_34_data_FIFO_blk[0] | proc_34_data_PIPO_blk[0] | proc_34_start_FIFO_blk[0] | proc_34_TLF_FIFO_blk[0] | proc_34_input_sync_blk[0] | proc_34_output_sync_blk[0]);
    assign proc_34_data_FIFO_blk[1] = 1'b0 | (~write_back63_U0.value_stream_V_V15_blk_n);
    assign proc_34_data_PIPO_blk[1] = 1'b0;
    assign proc_34_start_FIFO_blk[1] = 1'b0;
    assign proc_34_TLF_FIFO_blk[1] = 1'b0;
    assign proc_34_input_sync_blk[1] = 1'b0;
    assign proc_34_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_34[1] = dl_detect_out ? proc_dep_vld_vec_34_reg[1] : (proc_34_data_FIFO_blk[1] | proc_34_data_PIPO_blk[1] | proc_34_start_FIFO_blk[1] | proc_34_TLF_FIFO_blk[1] | proc_34_input_sync_blk[1] | proc_34_output_sync_blk[1]);
    assign proc_34_data_FIFO_blk[2] = 1'b0;
    assign proc_34_data_PIPO_blk[2] = 1'b0;
    assign proc_34_start_FIFO_blk[2] = 1'b0;
    assign proc_34_TLF_FIFO_blk[2] = 1'b0;
    assign proc_34_input_sync_blk[2] = 1'b0;
    assign proc_34_output_sync_blk[2] = 1'b0 | (ap_done_reg_15 & write_back63_U0.ap_done & ~write_back48_U0.ap_done);
    assign proc_dep_vld_vec_34[2] = dl_detect_out ? proc_dep_vld_vec_34_reg[2] : (proc_34_data_FIFO_blk[2] | proc_34_data_PIPO_blk[2] | proc_34_start_FIFO_blk[2] | proc_34_TLF_FIFO_blk[2] | proc_34_input_sync_blk[2] | proc_34_output_sync_blk[2]);
    assign proc_34_data_FIFO_blk[3] = 1'b0;
    assign proc_34_data_PIPO_blk[3] = 1'b0;
    assign proc_34_start_FIFO_blk[3] = 1'b0;
    assign proc_34_TLF_FIFO_blk[3] = 1'b0;
    assign proc_34_input_sync_blk[3] = 1'b0;
    assign proc_34_output_sync_blk[3] = 1'b0 | (ap_done_reg_15 & write_back63_U0.ap_done & ~write_back49_U0.ap_done);
    assign proc_dep_vld_vec_34[3] = dl_detect_out ? proc_dep_vld_vec_34_reg[3] : (proc_34_data_FIFO_blk[3] | proc_34_data_PIPO_blk[3] | proc_34_start_FIFO_blk[3] | proc_34_TLF_FIFO_blk[3] | proc_34_input_sync_blk[3] | proc_34_output_sync_blk[3]);
    assign proc_34_data_FIFO_blk[4] = 1'b0;
    assign proc_34_data_PIPO_blk[4] = 1'b0;
    assign proc_34_start_FIFO_blk[4] = 1'b0;
    assign proc_34_TLF_FIFO_blk[4] = 1'b0;
    assign proc_34_input_sync_blk[4] = 1'b0;
    assign proc_34_output_sync_blk[4] = 1'b0 | (ap_done_reg_15 & write_back63_U0.ap_done & ~write_back50_U0.ap_done);
    assign proc_dep_vld_vec_34[4] = dl_detect_out ? proc_dep_vld_vec_34_reg[4] : (proc_34_data_FIFO_blk[4] | proc_34_data_PIPO_blk[4] | proc_34_start_FIFO_blk[4] | proc_34_TLF_FIFO_blk[4] | proc_34_input_sync_blk[4] | proc_34_output_sync_blk[4]);
    assign proc_34_data_FIFO_blk[5] = 1'b0;
    assign proc_34_data_PIPO_blk[5] = 1'b0;
    assign proc_34_start_FIFO_blk[5] = 1'b0;
    assign proc_34_TLF_FIFO_blk[5] = 1'b0;
    assign proc_34_input_sync_blk[5] = 1'b0;
    assign proc_34_output_sync_blk[5] = 1'b0 | (ap_done_reg_15 & write_back63_U0.ap_done & ~write_back51_U0.ap_done);
    assign proc_dep_vld_vec_34[5] = dl_detect_out ? proc_dep_vld_vec_34_reg[5] : (proc_34_data_FIFO_blk[5] | proc_34_data_PIPO_blk[5] | proc_34_start_FIFO_blk[5] | proc_34_TLF_FIFO_blk[5] | proc_34_input_sync_blk[5] | proc_34_output_sync_blk[5]);
    assign proc_34_data_FIFO_blk[6] = 1'b0;
    assign proc_34_data_PIPO_blk[6] = 1'b0;
    assign proc_34_start_FIFO_blk[6] = 1'b0;
    assign proc_34_TLF_FIFO_blk[6] = 1'b0;
    assign proc_34_input_sync_blk[6] = 1'b0;
    assign proc_34_output_sync_blk[6] = 1'b0 | (ap_done_reg_15 & write_back63_U0.ap_done & ~write_back52_U0.ap_done);
    assign proc_dep_vld_vec_34[6] = dl_detect_out ? proc_dep_vld_vec_34_reg[6] : (proc_34_data_FIFO_blk[6] | proc_34_data_PIPO_blk[6] | proc_34_start_FIFO_blk[6] | proc_34_TLF_FIFO_blk[6] | proc_34_input_sync_blk[6] | proc_34_output_sync_blk[6]);
    assign proc_34_data_FIFO_blk[7] = 1'b0;
    assign proc_34_data_PIPO_blk[7] = 1'b0;
    assign proc_34_start_FIFO_blk[7] = 1'b0;
    assign proc_34_TLF_FIFO_blk[7] = 1'b0;
    assign proc_34_input_sync_blk[7] = 1'b0;
    assign proc_34_output_sync_blk[7] = 1'b0 | (ap_done_reg_15 & write_back63_U0.ap_done & ~write_back53_U0.ap_done);
    assign proc_dep_vld_vec_34[7] = dl_detect_out ? proc_dep_vld_vec_34_reg[7] : (proc_34_data_FIFO_blk[7] | proc_34_data_PIPO_blk[7] | proc_34_start_FIFO_blk[7] | proc_34_TLF_FIFO_blk[7] | proc_34_input_sync_blk[7] | proc_34_output_sync_blk[7]);
    assign proc_34_data_FIFO_blk[8] = 1'b0;
    assign proc_34_data_PIPO_blk[8] = 1'b0;
    assign proc_34_start_FIFO_blk[8] = 1'b0;
    assign proc_34_TLF_FIFO_blk[8] = 1'b0;
    assign proc_34_input_sync_blk[8] = 1'b0;
    assign proc_34_output_sync_blk[8] = 1'b0 | (ap_done_reg_15 & write_back63_U0.ap_done & ~write_back54_U0.ap_done);
    assign proc_dep_vld_vec_34[8] = dl_detect_out ? proc_dep_vld_vec_34_reg[8] : (proc_34_data_FIFO_blk[8] | proc_34_data_PIPO_blk[8] | proc_34_start_FIFO_blk[8] | proc_34_TLF_FIFO_blk[8] | proc_34_input_sync_blk[8] | proc_34_output_sync_blk[8]);
    assign proc_34_data_FIFO_blk[9] = 1'b0;
    assign proc_34_data_PIPO_blk[9] = 1'b0;
    assign proc_34_start_FIFO_blk[9] = 1'b0;
    assign proc_34_TLF_FIFO_blk[9] = 1'b0;
    assign proc_34_input_sync_blk[9] = 1'b0;
    assign proc_34_output_sync_blk[9] = 1'b0 | (ap_done_reg_15 & write_back63_U0.ap_done & ~write_back55_U0.ap_done);
    assign proc_dep_vld_vec_34[9] = dl_detect_out ? proc_dep_vld_vec_34_reg[9] : (proc_34_data_FIFO_blk[9] | proc_34_data_PIPO_blk[9] | proc_34_start_FIFO_blk[9] | proc_34_TLF_FIFO_blk[9] | proc_34_input_sync_blk[9] | proc_34_output_sync_blk[9]);
    assign proc_34_data_FIFO_blk[10] = 1'b0;
    assign proc_34_data_PIPO_blk[10] = 1'b0;
    assign proc_34_start_FIFO_blk[10] = 1'b0;
    assign proc_34_TLF_FIFO_blk[10] = 1'b0;
    assign proc_34_input_sync_blk[10] = 1'b0;
    assign proc_34_output_sync_blk[10] = 1'b0 | (ap_done_reg_15 & write_back63_U0.ap_done & ~write_back56_U0.ap_done);
    assign proc_dep_vld_vec_34[10] = dl_detect_out ? proc_dep_vld_vec_34_reg[10] : (proc_34_data_FIFO_blk[10] | proc_34_data_PIPO_blk[10] | proc_34_start_FIFO_blk[10] | proc_34_TLF_FIFO_blk[10] | proc_34_input_sync_blk[10] | proc_34_output_sync_blk[10]);
    assign proc_34_data_FIFO_blk[11] = 1'b0;
    assign proc_34_data_PIPO_blk[11] = 1'b0;
    assign proc_34_start_FIFO_blk[11] = 1'b0;
    assign proc_34_TLF_FIFO_blk[11] = 1'b0;
    assign proc_34_input_sync_blk[11] = 1'b0;
    assign proc_34_output_sync_blk[11] = 1'b0 | (ap_done_reg_15 & write_back63_U0.ap_done & ~write_back57_U0.ap_done);
    assign proc_dep_vld_vec_34[11] = dl_detect_out ? proc_dep_vld_vec_34_reg[11] : (proc_34_data_FIFO_blk[11] | proc_34_data_PIPO_blk[11] | proc_34_start_FIFO_blk[11] | proc_34_TLF_FIFO_blk[11] | proc_34_input_sync_blk[11] | proc_34_output_sync_blk[11]);
    assign proc_34_data_FIFO_blk[12] = 1'b0;
    assign proc_34_data_PIPO_blk[12] = 1'b0;
    assign proc_34_start_FIFO_blk[12] = 1'b0;
    assign proc_34_TLF_FIFO_blk[12] = 1'b0;
    assign proc_34_input_sync_blk[12] = 1'b0;
    assign proc_34_output_sync_blk[12] = 1'b0 | (ap_done_reg_15 & write_back63_U0.ap_done & ~write_back58_U0.ap_done);
    assign proc_dep_vld_vec_34[12] = dl_detect_out ? proc_dep_vld_vec_34_reg[12] : (proc_34_data_FIFO_blk[12] | proc_34_data_PIPO_blk[12] | proc_34_start_FIFO_blk[12] | proc_34_TLF_FIFO_blk[12] | proc_34_input_sync_blk[12] | proc_34_output_sync_blk[12]);
    assign proc_34_data_FIFO_blk[13] = 1'b0;
    assign proc_34_data_PIPO_blk[13] = 1'b0;
    assign proc_34_start_FIFO_blk[13] = 1'b0;
    assign proc_34_TLF_FIFO_blk[13] = 1'b0;
    assign proc_34_input_sync_blk[13] = 1'b0;
    assign proc_34_output_sync_blk[13] = 1'b0 | (ap_done_reg_15 & write_back63_U0.ap_done & ~write_back59_U0.ap_done);
    assign proc_dep_vld_vec_34[13] = dl_detect_out ? proc_dep_vld_vec_34_reg[13] : (proc_34_data_FIFO_blk[13] | proc_34_data_PIPO_blk[13] | proc_34_start_FIFO_blk[13] | proc_34_TLF_FIFO_blk[13] | proc_34_input_sync_blk[13] | proc_34_output_sync_blk[13]);
    assign proc_34_data_FIFO_blk[14] = 1'b0;
    assign proc_34_data_PIPO_blk[14] = 1'b0;
    assign proc_34_start_FIFO_blk[14] = 1'b0;
    assign proc_34_TLF_FIFO_blk[14] = 1'b0;
    assign proc_34_input_sync_blk[14] = 1'b0;
    assign proc_34_output_sync_blk[14] = 1'b0 | (ap_done_reg_15 & write_back63_U0.ap_done & ~write_back60_U0.ap_done);
    assign proc_dep_vld_vec_34[14] = dl_detect_out ? proc_dep_vld_vec_34_reg[14] : (proc_34_data_FIFO_blk[14] | proc_34_data_PIPO_blk[14] | proc_34_start_FIFO_blk[14] | proc_34_TLF_FIFO_blk[14] | proc_34_input_sync_blk[14] | proc_34_output_sync_blk[14]);
    assign proc_34_data_FIFO_blk[15] = 1'b0;
    assign proc_34_data_PIPO_blk[15] = 1'b0;
    assign proc_34_start_FIFO_blk[15] = 1'b0;
    assign proc_34_TLF_FIFO_blk[15] = 1'b0;
    assign proc_34_input_sync_blk[15] = 1'b0;
    assign proc_34_output_sync_blk[15] = 1'b0 | (ap_done_reg_15 & write_back63_U0.ap_done & ~write_back61_U0.ap_done);
    assign proc_dep_vld_vec_34[15] = dl_detect_out ? proc_dep_vld_vec_34_reg[15] : (proc_34_data_FIFO_blk[15] | proc_34_data_PIPO_blk[15] | proc_34_start_FIFO_blk[15] | proc_34_TLF_FIFO_blk[15] | proc_34_input_sync_blk[15] | proc_34_output_sync_blk[15]);
    assign proc_34_data_FIFO_blk[16] = 1'b0;
    assign proc_34_data_PIPO_blk[16] = 1'b0;
    assign proc_34_start_FIFO_blk[16] = 1'b0;
    assign proc_34_TLF_FIFO_blk[16] = 1'b0;
    assign proc_34_input_sync_blk[16] = 1'b0;
    assign proc_34_output_sync_blk[16] = 1'b0 | (ap_done_reg_15 & write_back63_U0.ap_done & ~write_back62_U0.ap_done);
    assign proc_dep_vld_vec_34[16] = dl_detect_out ? proc_dep_vld_vec_34_reg[16] : (proc_34_data_FIFO_blk[16] | proc_34_data_PIPO_blk[16] | proc_34_start_FIFO_blk[16] | proc_34_TLF_FIFO_blk[16] | proc_34_input_sync_blk[16] | proc_34_output_sync_blk[16]);
    always @ (negedge reset or posedge clock) begin
        if (~reset) begin
            proc_dep_vld_vec_34_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_34_reg <= proc_dep_vld_vec_34;
        end
    end
    assign in_chan_dep_vld_vec_34[0] = dep_chan_vld_0_34;
    assign in_chan_dep_data_vec_34[34 : 0] = dep_chan_data_0_34;
    assign token_in_vec_34[0] = token_0_34;
    assign in_chan_dep_vld_vec_34[1] = dep_chan_vld_18_34;
    assign in_chan_dep_data_vec_34[69 : 35] = dep_chan_data_18_34;
    assign token_in_vec_34[1] = token_18_34;
    assign in_chan_dep_vld_vec_34[2] = dep_chan_vld_19_34;
    assign in_chan_dep_data_vec_34[104 : 70] = dep_chan_data_19_34;
    assign token_in_vec_34[2] = token_19_34;
    assign in_chan_dep_vld_vec_34[3] = dep_chan_vld_20_34;
    assign in_chan_dep_data_vec_34[139 : 105] = dep_chan_data_20_34;
    assign token_in_vec_34[3] = token_20_34;
    assign in_chan_dep_vld_vec_34[4] = dep_chan_vld_21_34;
    assign in_chan_dep_data_vec_34[174 : 140] = dep_chan_data_21_34;
    assign token_in_vec_34[4] = token_21_34;
    assign in_chan_dep_vld_vec_34[5] = dep_chan_vld_22_34;
    assign in_chan_dep_data_vec_34[209 : 175] = dep_chan_data_22_34;
    assign token_in_vec_34[5] = token_22_34;
    assign in_chan_dep_vld_vec_34[6] = dep_chan_vld_23_34;
    assign in_chan_dep_data_vec_34[244 : 210] = dep_chan_data_23_34;
    assign token_in_vec_34[6] = token_23_34;
    assign in_chan_dep_vld_vec_34[7] = dep_chan_vld_24_34;
    assign in_chan_dep_data_vec_34[279 : 245] = dep_chan_data_24_34;
    assign token_in_vec_34[7] = token_24_34;
    assign in_chan_dep_vld_vec_34[8] = dep_chan_vld_25_34;
    assign in_chan_dep_data_vec_34[314 : 280] = dep_chan_data_25_34;
    assign token_in_vec_34[8] = token_25_34;
    assign in_chan_dep_vld_vec_34[9] = dep_chan_vld_26_34;
    assign in_chan_dep_data_vec_34[349 : 315] = dep_chan_data_26_34;
    assign token_in_vec_34[9] = token_26_34;
    assign in_chan_dep_vld_vec_34[10] = dep_chan_vld_27_34;
    assign in_chan_dep_data_vec_34[384 : 350] = dep_chan_data_27_34;
    assign token_in_vec_34[10] = token_27_34;
    assign in_chan_dep_vld_vec_34[11] = dep_chan_vld_28_34;
    assign in_chan_dep_data_vec_34[419 : 385] = dep_chan_data_28_34;
    assign token_in_vec_34[11] = token_28_34;
    assign in_chan_dep_vld_vec_34[12] = dep_chan_vld_29_34;
    assign in_chan_dep_data_vec_34[454 : 420] = dep_chan_data_29_34;
    assign token_in_vec_34[12] = token_29_34;
    assign in_chan_dep_vld_vec_34[13] = dep_chan_vld_30_34;
    assign in_chan_dep_data_vec_34[489 : 455] = dep_chan_data_30_34;
    assign token_in_vec_34[13] = token_30_34;
    assign in_chan_dep_vld_vec_34[14] = dep_chan_vld_31_34;
    assign in_chan_dep_data_vec_34[524 : 490] = dep_chan_data_31_34;
    assign token_in_vec_34[14] = token_31_34;
    assign in_chan_dep_vld_vec_34[15] = dep_chan_vld_32_34;
    assign in_chan_dep_data_vec_34[559 : 525] = dep_chan_data_32_34;
    assign token_in_vec_34[15] = token_32_34;
    assign in_chan_dep_vld_vec_34[16] = dep_chan_vld_33_34;
    assign in_chan_dep_data_vec_34[594 : 560] = dep_chan_data_33_34;
    assign token_in_vec_34[16] = token_33_34;
    assign dep_chan_vld_34_0 = out_chan_dep_vld_vec_34[0];
    assign dep_chan_data_34_0 = out_chan_dep_data_34;
    assign token_34_0 = token_out_vec_34[0];
    assign dep_chan_vld_34_18 = out_chan_dep_vld_vec_34[1];
    assign dep_chan_data_34_18 = out_chan_dep_data_34;
    assign token_34_18 = token_out_vec_34[1];
    assign dep_chan_vld_34_19 = out_chan_dep_vld_vec_34[2];
    assign dep_chan_data_34_19 = out_chan_dep_data_34;
    assign token_34_19 = token_out_vec_34[2];
    assign dep_chan_vld_34_20 = out_chan_dep_vld_vec_34[3];
    assign dep_chan_data_34_20 = out_chan_dep_data_34;
    assign token_34_20 = token_out_vec_34[3];
    assign dep_chan_vld_34_21 = out_chan_dep_vld_vec_34[4];
    assign dep_chan_data_34_21 = out_chan_dep_data_34;
    assign token_34_21 = token_out_vec_34[4];
    assign dep_chan_vld_34_22 = out_chan_dep_vld_vec_34[5];
    assign dep_chan_data_34_22 = out_chan_dep_data_34;
    assign token_34_22 = token_out_vec_34[5];
    assign dep_chan_vld_34_23 = out_chan_dep_vld_vec_34[6];
    assign dep_chan_data_34_23 = out_chan_dep_data_34;
    assign token_34_23 = token_out_vec_34[6];
    assign dep_chan_vld_34_24 = out_chan_dep_vld_vec_34[7];
    assign dep_chan_data_34_24 = out_chan_dep_data_34;
    assign token_34_24 = token_out_vec_34[7];
    assign dep_chan_vld_34_25 = out_chan_dep_vld_vec_34[8];
    assign dep_chan_data_34_25 = out_chan_dep_data_34;
    assign token_34_25 = token_out_vec_34[8];
    assign dep_chan_vld_34_26 = out_chan_dep_vld_vec_34[9];
    assign dep_chan_data_34_26 = out_chan_dep_data_34;
    assign token_34_26 = token_out_vec_34[9];
    assign dep_chan_vld_34_27 = out_chan_dep_vld_vec_34[10];
    assign dep_chan_data_34_27 = out_chan_dep_data_34;
    assign token_34_27 = token_out_vec_34[10];
    assign dep_chan_vld_34_28 = out_chan_dep_vld_vec_34[11];
    assign dep_chan_data_34_28 = out_chan_dep_data_34;
    assign token_34_28 = token_out_vec_34[11];
    assign dep_chan_vld_34_29 = out_chan_dep_vld_vec_34[12];
    assign dep_chan_data_34_29 = out_chan_dep_data_34;
    assign token_34_29 = token_out_vec_34[12];
    assign dep_chan_vld_34_30 = out_chan_dep_vld_vec_34[13];
    assign dep_chan_data_34_30 = out_chan_dep_data_34;
    assign token_34_30 = token_out_vec_34[13];
    assign dep_chan_vld_34_31 = out_chan_dep_vld_vec_34[14];
    assign dep_chan_data_34_31 = out_chan_dep_data_34;
    assign token_34_31 = token_out_vec_34[14];
    assign dep_chan_vld_34_32 = out_chan_dep_vld_vec_34[15];
    assign dep_chan_data_34_32 = out_chan_dep_data_34;
    assign token_34_32 = token_out_vec_34[15];
    assign dep_chan_vld_34_33 = out_chan_dep_vld_vec_34[16];
    assign dep_chan_data_34_33 = out_chan_dep_data_34;
    assign token_34_33 = token_out_vec_34[16];


`include "kernel_pr_hls_deadlock_report_unit.vh"
